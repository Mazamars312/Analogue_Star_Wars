`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.05.2023 09:26:30
// Design Name: 
// Module Name: Sound_program_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sound_program_rom_1(
    input               clk,
    input       [13:0]  address,
    output reg  [7:0]   data
    );
    
    reg [7:0] ROM_MEM [16383:0];
    
    integer i;
    initial begin
        ROM_MEM[0   ] = 8'hBE;
ROM_MEM[1   ] = 8'hE4;
ROM_MEM[2   ] = 8'h40;
ROM_MEM[3   ] = 8'h62;
ROM_MEM[4   ] = 8'h41;
ROM_MEM[5   ] = 8'h9B;
ROM_MEM[6   ] = 8'h40;
ROM_MEM[7   ] = 8'h62;
ROM_MEM[8   ] = 8'h41;
ROM_MEM[9   ] = 8'h9B;
ROM_MEM[10  ] = 8'h41;
ROM_MEM[11  ] = 8'h9C;
ROM_MEM[12  ] = 8'h42;
ROM_MEM[13  ] = 8'h40;
ROM_MEM[14  ] = 8'h42;
ROM_MEM[15  ] = 8'h41;
ROM_MEM[16  ] = 8'h42;
ROM_MEM[17  ] = 8'hFB;
ROM_MEM[18  ] = 8'h42;
ROM_MEM[19  ] = 8'hFC;
ROM_MEM[20  ] = 8'h44;
ROM_MEM[21  ] = 8'h35;
ROM_MEM[22  ] = 8'h44;
ROM_MEM[23  ] = 8'h36;
ROM_MEM[24  ] = 8'h45;
ROM_MEM[25  ] = 8'h76;
ROM_MEM[26  ] = 8'h45;
ROM_MEM[27  ] = 8'h77;
ROM_MEM[28  ] = 8'h46;
ROM_MEM[29  ] = 8'hC2;
ROM_MEM[30  ] = 8'h46;
ROM_MEM[31  ] = 8'hC3;
ROM_MEM[32  ] = 8'h48;
ROM_MEM[33  ] = 8'h02;
ROM_MEM[34  ] = 8'h48;
ROM_MEM[35  ] = 8'h03;
ROM_MEM[36  ] = 8'h48;
ROM_MEM[37  ] = 8'hDF;
ROM_MEM[38  ] = 8'h48;
ROM_MEM[39  ] = 8'hE0;
ROM_MEM[40  ] = 8'h49;
ROM_MEM[41  ] = 8'hD5;
ROM_MEM[42  ] = 8'h49;
ROM_MEM[43  ] = 8'hD6;
ROM_MEM[44  ] = 8'h4A;
ROM_MEM[45  ] = 8'h58;
ROM_MEM[46  ] = 8'h4A;
ROM_MEM[47  ] = 8'h59;
ROM_MEM[48  ] = 8'h4B;
ROM_MEM[49  ] = 8'h37;
ROM_MEM[50  ] = 8'h4B;
ROM_MEM[51  ] = 8'h38;
ROM_MEM[52  ] = 8'h4C;
ROM_MEM[53  ] = 8'h49;
ROM_MEM[54  ] = 8'h4C;
ROM_MEM[55  ] = 8'h4A;
ROM_MEM[56  ] = 8'h4D;
ROM_MEM[57  ] = 8'hB9;
ROM_MEM[58  ] = 8'h4D;
ROM_MEM[59  ] = 8'hBA;
ROM_MEM[60  ] = 8'h4F;
ROM_MEM[61  ] = 8'h30;
ROM_MEM[62  ] = 8'h4F;
ROM_MEM[63  ] = 8'h31;
ROM_MEM[64  ] = 8'h50;
ROM_MEM[65  ] = 8'h2D;
ROM_MEM[66  ] = 8'h50;
ROM_MEM[67  ] = 8'h2E;
ROM_MEM[68  ] = 8'h50;
ROM_MEM[69  ] = 8'hA6;
ROM_MEM[70  ] = 8'h50;
ROM_MEM[71  ] = 8'hA7;
ROM_MEM[72  ] = 8'h51;
ROM_MEM[73  ] = 8'hA3;
ROM_MEM[74  ] = 8'h51;
ROM_MEM[75  ] = 8'hA4;
ROM_MEM[76  ] = 8'h52;
ROM_MEM[77  ] = 8'hC7;
ROM_MEM[78  ] = 8'h52;
ROM_MEM[79  ] = 8'hC8;
ROM_MEM[80  ] = 8'h54;
ROM_MEM[81  ] = 8'hC8;
ROM_MEM[82  ] = 8'h54;
ROM_MEM[83  ] = 8'hCD;
ROM_MEM[84  ] = 8'h55;
ROM_MEM[85  ] = 8'h7C;
ROM_MEM[86  ] = 8'h55;
ROM_MEM[87  ] = 8'h7D;
ROM_MEM[88  ] = 8'h57;
ROM_MEM[89  ] = 8'h46;
ROM_MEM[90  ] = 8'h57;
ROM_MEM[91  ] = 8'h47;
ROM_MEM[92  ] = 8'h58;
ROM_MEM[93  ] = 8'h0F;
ROM_MEM[94  ] = 8'h58;
ROM_MEM[95  ] = 8'h10;
ROM_MEM[96  ] = 8'h58;
ROM_MEM[97  ] = 8'hE4;
ROM_MEM[98  ] = 8'h04;
ROM_MEM[99  ] = 8'h00;
ROM_MEM[100 ] = 8'h7A;
ROM_MEM[101 ] = 8'h8A;
ROM_MEM[102 ] = 8'h01;
ROM_MEM[103 ] = 8'hC0;
ROM_MEM[104 ] = 8'h4F;
ROM_MEM[105 ] = 8'h33;
ROM_MEM[106 ] = 8'h80;
ROM_MEM[107 ] = 8'h68;
ROM_MEM[108 ] = 8'h99;
ROM_MEM[109 ] = 8'h50;
ROM_MEM[110 ] = 8'h67;
ROM_MEM[111 ] = 8'h8D;
ROM_MEM[112 ] = 8'h9E;
ROM_MEM[113 ] = 8'h95;
ROM_MEM[114 ] = 8'hB5;
ROM_MEM[115 ] = 8'h5A;
ROM_MEM[116 ] = 8'h9E;
ROM_MEM[117 ] = 8'h8D;
ROM_MEM[118 ] = 8'hA8;
ROM_MEM[119 ] = 8'h86;
ROM_MEM[120 ] = 8'h4F;
ROM_MEM[121 ] = 8'h6E;
ROM_MEM[122 ] = 8'h49;
ROM_MEM[123 ] = 8'h34;
ROM_MEM[124 ] = 8'hEE;
ROM_MEM[125 ] = 8'h6A;
ROM_MEM[126 ] = 8'hD1;
ROM_MEM[127 ] = 8'hA8;
ROM_MEM[128 ] = 8'h44;
ROM_MEM[129 ] = 8'hC1;
ROM_MEM[130 ] = 8'h44;
ROM_MEM[131 ] = 8'hB2;
ROM_MEM[132 ] = 8'hF8;
ROM_MEM[133 ] = 8'h92;
ROM_MEM[134 ] = 8'h12;
ROM_MEM[135 ] = 8'h78;
ROM_MEM[136 ] = 8'h5F;
ROM_MEM[137 ] = 8'h41;
ROM_MEM[138 ] = 8'h6A;
ROM_MEM[139 ] = 8'h4B;
ROM_MEM[140 ] = 8'h8B;
ROM_MEM[141 ] = 8'hEF;
ROM_MEM[142 ] = 8'h7D;
ROM_MEM[143 ] = 8'h27;
ROM_MEM[144 ] = 8'h89;
ROM_MEM[145 ] = 8'hCD;
ROM_MEM[146 ] = 8'h2B;
ROM_MEM[147 ] = 8'hBE;
ROM_MEM[148 ] = 8'h8F;
ROM_MEM[149 ] = 8'h95;
ROM_MEM[150 ] = 8'hA8;
ROM_MEM[151 ] = 8'hD6;
ROM_MEM[152 ] = 8'hAE;
ROM_MEM[153 ] = 8'hF8;
ROM_MEM[154 ] = 8'hDE;
ROM_MEM[155 ] = 8'h57;
ROM_MEM[156 ] = 8'h81;
ROM_MEM[157 ] = 8'hD8;
ROM_MEM[158 ] = 8'hBA;
ROM_MEM[159 ] = 8'hE2;
ROM_MEM[160 ] = 8'h07;
ROM_MEM[161 ] = 8'h13;
ROM_MEM[162 ] = 8'h43;
ROM_MEM[163 ] = 8'hA2;
ROM_MEM[164 ] = 8'hED;
ROM_MEM[165 ] = 8'h8A;
ROM_MEM[166 ] = 8'h1F;
ROM_MEM[167 ] = 8'hA5;
ROM_MEM[168 ] = 8'h36;
ROM_MEM[169 ] = 8'hBB;
ROM_MEM[170 ] = 8'hAE;
ROM_MEM[171 ] = 8'h2A;
ROM_MEM[172 ] = 8'h41;
ROM_MEM[173 ] = 8'h34;
ROM_MEM[174 ] = 8'h66;
ROM_MEM[175 ] = 8'h92;
ROM_MEM[176 ] = 8'hD1;
ROM_MEM[177 ] = 8'hB8;
ROM_MEM[178 ] = 8'h24;
ROM_MEM[179 ] = 8'h55;
ROM_MEM[180 ] = 8'hBB;
ROM_MEM[181 ] = 8'h09;
ROM_MEM[182 ] = 8'h5B;
ROM_MEM[183 ] = 8'h92;
ROM_MEM[184 ] = 8'h92;
ROM_MEM[185 ] = 8'h4F;
ROM_MEM[186 ] = 8'h67;
ROM_MEM[187 ] = 8'h6A;
ROM_MEM[188 ] = 8'hAC;
ROM_MEM[189 ] = 8'h56;
ROM_MEM[190 ] = 8'h0C;
ROM_MEM[191 ] = 8'h10;
ROM_MEM[192 ] = 8'h29;
ROM_MEM[193 ] = 8'h8B;
ROM_MEM[194 ] = 8'h01;
ROM_MEM[195 ] = 8'h0A;
ROM_MEM[196 ] = 8'h46;
ROM_MEM[197 ] = 8'h35;
ROM_MEM[198 ] = 8'h40;
ROM_MEM[199 ] = 8'h82;
ROM_MEM[200 ] = 8'h6C;
ROM_MEM[201 ] = 8'h0A;
ROM_MEM[202 ] = 8'h08;
ROM_MEM[203 ] = 8'h50;
ROM_MEM[204 ] = 8'h98;
ROM_MEM[205 ] = 8'h01;
ROM_MEM[206 ] = 8'h1C;
ROM_MEM[207 ] = 8'hB2;
ROM_MEM[208 ] = 8'h2A;
ROM_MEM[209 ] = 8'h80;
ROM_MEM[210 ] = 8'hD0;
ROM_MEM[211 ] = 8'hCA;
ROM_MEM[212 ] = 8'h54;
ROM_MEM[213 ] = 8'h66;
ROM_MEM[214 ] = 8'h95;
ROM_MEM[215 ] = 8'h49;
ROM_MEM[216 ] = 8'h32;
ROM_MEM[217 ] = 8'h91;
ROM_MEM[218 ] = 8'h73;
ROM_MEM[219 ] = 8'hA9;
ROM_MEM[220 ] = 8'h00;
ROM_MEM[221 ] = 8'h11;
ROM_MEM[222 ] = 8'h5C;
ROM_MEM[223 ] = 8'h18;
ROM_MEM[224 ] = 8'h00;
ROM_MEM[225 ] = 8'h64;
ROM_MEM[226 ] = 8'h06;
ROM_MEM[227 ] = 8'h01;
ROM_MEM[228 ] = 8'h80;
ROM_MEM[229 ] = 8'h50;
ROM_MEM[230 ] = 8'h65;
ROM_MEM[231 ] = 8'h00;
ROM_MEM[232 ] = 8'h61;
ROM_MEM[233 ] = 8'h2A;
ROM_MEM[234 ] = 8'h02;
ROM_MEM[235 ] = 8'h60;
ROM_MEM[236 ] = 8'h42;
ROM_MEM[237 ] = 8'h55;
ROM_MEM[238 ] = 8'h00;
ROM_MEM[239 ] = 8'h4C;
ROM_MEM[240 ] = 8'h99;
ROM_MEM[241 ] = 8'h86;
ROM_MEM[242 ] = 8'h2C;
ROM_MEM[243 ] = 8'hF8;
ROM_MEM[244 ] = 8'h29;
ROM_MEM[245 ] = 8'h66;
ROM_MEM[246 ] = 8'hAB;
ROM_MEM[247 ] = 8'hDD;
ROM_MEM[248 ] = 8'h92;
ROM_MEM[249 ] = 8'hE8;
ROM_MEM[250 ] = 8'h76;
ROM_MEM[251 ] = 8'h84;
ROM_MEM[252 ] = 8'hA5;
ROM_MEM[253 ] = 8'h4A;
ROM_MEM[254 ] = 8'h8B;
ROM_MEM[255 ] = 8'h92;
ROM_MEM[256 ] = 8'hDE;
ROM_MEM[257 ] = 8'h11;
ROM_MEM[258 ] = 8'hE6;
ROM_MEM[259 ] = 8'h29;
ROM_MEM[260 ] = 8'h23;
ROM_MEM[261 ] = 8'h88;
ROM_MEM[262 ] = 8'h66;
ROM_MEM[263 ] = 8'h47;
ROM_MEM[264 ] = 8'h54;
ROM_MEM[265 ] = 8'hA7;
ROM_MEM[266 ] = 8'h0C;
ROM_MEM[267 ] = 8'h3F;
ROM_MEM[268 ] = 8'hA4;
ROM_MEM[269 ] = 8'h6B;
ROM_MEM[270 ] = 8'h71;
ROM_MEM[271 ] = 8'hAD;
ROM_MEM[272 ] = 8'h37;
ROM_MEM[273 ] = 8'hFC;
ROM_MEM[274 ] = 8'h10;
ROM_MEM[275 ] = 8'h77;
ROM_MEM[276 ] = 8'h44;
ROM_MEM[277 ] = 8'hBD;
ROM_MEM[278 ] = 8'h5A;
ROM_MEM[279 ] = 8'hF3;
ROM_MEM[280 ] = 8'hA3;
ROM_MEM[281 ] = 8'hDB;
ROM_MEM[282 ] = 8'h15;
ROM_MEM[283 ] = 8'hB3;
ROM_MEM[284 ] = 8'hAA;
ROM_MEM[285 ] = 8'h2D;
ROM_MEM[286 ] = 8'hC8;
ROM_MEM[287 ] = 8'hBA;
ROM_MEM[288 ] = 8'h96;
ROM_MEM[289 ] = 8'hD9;
ROM_MEM[290 ] = 8'h4A;
ROM_MEM[291 ] = 8'hA7;
ROM_MEM[292 ] = 8'h38;
ROM_MEM[293 ] = 8'hDA;
ROM_MEM[294 ] = 8'h1E;
ROM_MEM[295 ] = 8'h54;
ROM_MEM[296 ] = 8'h8F;
ROM_MEM[297 ] = 8'h2C;
ROM_MEM[298 ] = 8'h00;
ROM_MEM[299 ] = 8'h16;
ROM_MEM[300 ] = 8'h5D;
ROM_MEM[301 ] = 8'h18;
ROM_MEM[302 ] = 8'h40;
ROM_MEM[303 ] = 8'h49;
ROM_MEM[304 ] = 8'hA4;
ROM_MEM[305 ] = 8'h01;
ROM_MEM[306 ] = 8'h0A;
ROM_MEM[307 ] = 8'h24;
ROM_MEM[308 ] = 8'h73;
ROM_MEM[309 ] = 8'h40;
ROM_MEM[310 ] = 8'h81;
ROM_MEM[311 ] = 8'h62;
ROM_MEM[312 ] = 8'h06;
ROM_MEM[313 ] = 8'h48;
ROM_MEM[314 ] = 8'h40;
ROM_MEM[315 ] = 8'hD9;
ROM_MEM[316 ] = 8'h01;
ROM_MEM[317 ] = 8'h19;
ROM_MEM[318 ] = 8'hA9;
ROM_MEM[319 ] = 8'h38;
ROM_MEM[320 ] = 8'hA0;
ROM_MEM[321 ] = 8'h40;
ROM_MEM[322 ] = 8'h51;
ROM_MEM[323 ] = 8'h05;
ROM_MEM[324 ] = 8'h04;
ROM_MEM[325 ] = 8'hC8;
ROM_MEM[326 ] = 8'h42;
ROM_MEM[327 ] = 8'h00;
ROM_MEM[328 ] = 8'h00;
ROM_MEM[329 ] = 8'hD9;
ROM_MEM[330 ] = 8'h18;
ROM_MEM[331 ] = 8'h40;
ROM_MEM[332 ] = 8'hB1;
ROM_MEM[333 ] = 8'h25;
ROM_MEM[334 ] = 8'h03;
ROM_MEM[335 ] = 8'h80;
ROM_MEM[336 ] = 8'hA9;
ROM_MEM[337 ] = 8'h10;
ROM_MEM[338 ] = 8'h00;
ROM_MEM[339 ] = 8'h88;
ROM_MEM[340 ] = 8'h95;
ROM_MEM[341 ] = 8'hA9;
ROM_MEM[342 ] = 8'hCE;
ROM_MEM[343 ] = 8'h52;
ROM_MEM[344 ] = 8'h4A;
ROM_MEM[345 ] = 8'h3C;
ROM_MEM[346 ] = 8'h92;
ROM_MEM[347 ] = 8'h94;
ROM_MEM[348 ] = 8'h32;
ROM_MEM[349 ] = 8'h6A;
ROM_MEM[350 ] = 8'h2F;
ROM_MEM[351 ] = 8'h31;
ROM_MEM[352 ] = 8'h6F;
ROM_MEM[353 ] = 8'h94;
ROM_MEM[354 ] = 8'h52;
ROM_MEM[355 ] = 8'h67;
ROM_MEM[356 ] = 8'h2B;
ROM_MEM[357 ] = 8'h25;
ROM_MEM[358 ] = 8'hBC;
ROM_MEM[359 ] = 8'h49;
ROM_MEM[360 ] = 8'h09;
ROM_MEM[361 ] = 8'h83;
ROM_MEM[362 ] = 8'hF4;
ROM_MEM[363 ] = 8'h36;
ROM_MEM[364 ] = 8'hE5;
ROM_MEM[365 ] = 8'hA6;
ROM_MEM[366 ] = 8'hC5;
ROM_MEM[367 ] = 8'h77;
ROM_MEM[368 ] = 8'h36;
ROM_MEM[369 ] = 8'h4B;
ROM_MEM[370 ] = 8'h4D;
ROM_MEM[371 ] = 8'h9A;
ROM_MEM[372 ] = 8'h05;
ROM_MEM[373 ] = 8'hDF;
ROM_MEM[374 ] = 8'h84;
ROM_MEM[375 ] = 8'h2C;
ROM_MEM[376 ] = 8'h52;
ROM_MEM[377 ] = 8'h5B;
ROM_MEM[378 ] = 8'hEB;
ROM_MEM[379 ] = 8'hC2;
ROM_MEM[380 ] = 8'hE0;
ROM_MEM[381 ] = 8'hBB;
ROM_MEM[382 ] = 8'h4C;
ROM_MEM[383 ] = 8'h49;
ROM_MEM[384 ] = 8'h29;
ROM_MEM[385 ] = 8'h03;
ROM_MEM[386 ] = 8'h80;
ROM_MEM[387 ] = 8'h29;
ROM_MEM[388 ] = 8'h27;
ROM_MEM[389 ] = 8'h00;
ROM_MEM[390 ] = 8'hD0;
ROM_MEM[391 ] = 8'h1D;
ROM_MEM[392 ] = 8'h04;
ROM_MEM[393 ] = 8'h00;
ROM_MEM[394 ] = 8'hB2;
ROM_MEM[395 ] = 8'h13;
ROM_MEM[396 ] = 8'h80;
ROM_MEM[397 ] = 8'h01;
ROM_MEM[398 ] = 8'h3A;
ROM_MEM[399 ] = 8'h13;
ROM_MEM[400 ] = 8'h09;
ROM_MEM[401 ] = 8'h40;
ROM_MEM[402 ] = 8'h27;
ROM_MEM[403 ] = 8'h22;
ROM_MEM[404 ] = 8'h02;
ROM_MEM[405 ] = 8'h80;
ROM_MEM[406 ] = 8'h10;
ROM_MEM[407 ] = 8'hF2;
ROM_MEM[408 ] = 8'h00;
ROM_MEM[409 ] = 8'h50;
ROM_MEM[410 ] = 8'h58;
ROM_MEM[411 ] = 8'h01;
ROM_MEM[412 ] = 8'h04;
ROM_MEM[413 ] = 8'h00;
ROM_MEM[414 ] = 8'hA2;
ROM_MEM[415 ] = 8'h82;
ROM_MEM[416 ] = 8'h01;
ROM_MEM[417 ] = 8'h38;
ROM_MEM[418 ] = 8'hAB;
ROM_MEM[419 ] = 8'h30;
ROM_MEM[420 ] = 8'h80;
ROM_MEM[421 ] = 8'h65;
ROM_MEM[422 ] = 8'hB2;
ROM_MEM[423 ] = 8'hD0;
ROM_MEM[424 ] = 8'hA5;
ROM_MEM[425 ] = 8'hA1;
ROM_MEM[426 ] = 8'hEC;
ROM_MEM[427 ] = 8'h61;
ROM_MEM[428 ] = 8'h69;
ROM_MEM[429 ] = 8'h52;
ROM_MEM[430 ] = 8'h97;
ROM_MEM[431 ] = 8'h8A;
ROM_MEM[432 ] = 8'hBA;
ROM_MEM[433 ] = 8'hB1;
ROM_MEM[434 ] = 8'hB7;
ROM_MEM[435 ] = 8'h72;
ROM_MEM[436 ] = 8'h7D;
ROM_MEM[437 ] = 8'h50;
ROM_MEM[438 ] = 8'hA1;
ROM_MEM[439 ] = 8'h12;
ROM_MEM[440 ] = 8'h99;
ROM_MEM[441 ] = 8'hD6;
ROM_MEM[442 ] = 8'h35;
ROM_MEM[443 ] = 8'h8E;
ROM_MEM[444 ] = 8'h7B;
ROM_MEM[445 ] = 8'h44;
ROM_MEM[446 ] = 8'h7A;
ROM_MEM[447 ] = 8'h9A;
ROM_MEM[448 ] = 8'h50;
ROM_MEM[449 ] = 8'h39;
ROM_MEM[450 ] = 8'hE1;
ROM_MEM[451 ] = 8'h91;
ROM_MEM[452 ] = 8'h61;
ROM_MEM[453 ] = 8'h89;
ROM_MEM[454 ] = 8'h57;
ROM_MEM[455 ] = 8'h51;
ROM_MEM[456 ] = 8'h5D;
ROM_MEM[457 ] = 8'hBA;
ROM_MEM[458 ] = 8'h88;
ROM_MEM[459 ] = 8'h4D;
ROM_MEM[460 ] = 8'h3E;
ROM_MEM[461 ] = 8'h79;
ROM_MEM[462 ] = 8'hB3;
ROM_MEM[463 ] = 8'h19;
ROM_MEM[464 ] = 8'h2A;
ROM_MEM[465 ] = 8'h3E;
ROM_MEM[466 ] = 8'hFA;
ROM_MEM[467 ] = 8'hE4;
ROM_MEM[468 ] = 8'hCD;
ROM_MEM[469 ] = 8'h55;
ROM_MEM[470 ] = 8'h1A;
ROM_MEM[471 ] = 8'hD9;
ROM_MEM[472 ] = 8'hA4;
ROM_MEM[473 ] = 8'h93;
ROM_MEM[474 ] = 8'h35;
ROM_MEM[475 ] = 8'h9B;
ROM_MEM[476 ] = 8'h69;
ROM_MEM[477 ] = 8'h2C;
ROM_MEM[478 ] = 8'h93;
ROM_MEM[479 ] = 8'h5A;
ROM_MEM[480 ] = 8'h96;
ROM_MEM[481 ] = 8'h8C;
ROM_MEM[482 ] = 8'h19;
ROM_MEM[483 ] = 8'h6B;
ROM_MEM[484 ] = 8'h54;
ROM_MEM[485 ] = 8'h2D;
ROM_MEM[486 ] = 8'h99;
ROM_MEM[487 ] = 8'hD7;
ROM_MEM[488 ] = 8'hE6;
ROM_MEM[489 ] = 8'hEA;
ROM_MEM[490 ] = 8'h19;
ROM_MEM[491 ] = 8'hB7;
ROM_MEM[492 ] = 8'h64;
ROM_MEM[493 ] = 8'hCE;
ROM_MEM[494 ] = 8'h5A;
ROM_MEM[495 ] = 8'h88;
ROM_MEM[496 ] = 8'h46;
ROM_MEM[497 ] = 8'hB3;
ROM_MEM[498 ] = 8'h92;
ROM_MEM[499 ] = 8'h3B;
ROM_MEM[500 ] = 8'hEB;
ROM_MEM[501 ] = 8'h2E;
ROM_MEM[502 ] = 8'h1A;
ROM_MEM[503 ] = 8'hED;
ROM_MEM[504 ] = 8'h52;
ROM_MEM[505 ] = 8'h61;
ROM_MEM[506 ] = 8'hBC;
ROM_MEM[507 ] = 8'h9B;
ROM_MEM[508 ] = 8'hAA;
ROM_MEM[509 ] = 8'hB7;
ROM_MEM[510 ] = 8'h0D;
ROM_MEM[511 ] = 8'h95;
ROM_MEM[512 ] = 8'h33;
ROM_MEM[513 ] = 8'hE1;
ROM_MEM[514 ] = 8'hA2;
ROM_MEM[515 ] = 8'hD1;
ROM_MEM[516 ] = 8'h64;
ROM_MEM[517 ] = 8'h14;
ROM_MEM[518 ] = 8'hD9;
ROM_MEM[519 ] = 8'h66;
ROM_MEM[520 ] = 8'h08;
ROM_MEM[521 ] = 8'hDB;
ROM_MEM[522 ] = 8'hEC;
ROM_MEM[523 ] = 8'h55;
ROM_MEM[524 ] = 8'h16;
ROM_MEM[525 ] = 8'h93;
ROM_MEM[526 ] = 8'hA1;
ROM_MEM[527 ] = 8'h6C;
ROM_MEM[528 ] = 8'hB7;
ROM_MEM[529 ] = 8'h57;
ROM_MEM[530 ] = 8'h55;
ROM_MEM[531 ] = 8'h6C;
ROM_MEM[532 ] = 8'hBA;
ROM_MEM[533 ] = 8'h92;
ROM_MEM[534 ] = 8'h5F;
ROM_MEM[535 ] = 8'h59;
ROM_MEM[536 ] = 8'h55;
ROM_MEM[537 ] = 8'h71;
ROM_MEM[538 ] = 8'h15;
ROM_MEM[539 ] = 8'h4A;
ROM_MEM[540 ] = 8'h3E;
ROM_MEM[541 ] = 8'h65;
ROM_MEM[542 ] = 8'hD5;
ROM_MEM[543 ] = 8'hC5;
ROM_MEM[544 ] = 8'h97;
ROM_MEM[545 ] = 8'h2B;
ROM_MEM[546 ] = 8'hE7;
ROM_MEM[547 ] = 8'h94;
ROM_MEM[548 ] = 8'hD1;
ROM_MEM[549 ] = 8'hE4;
ROM_MEM[550 ] = 8'h10;
ROM_MEM[551 ] = 8'h29;
ROM_MEM[552 ] = 8'h32;
ROM_MEM[553 ] = 8'h55;
ROM_MEM[554 ] = 8'h46;
ROM_MEM[555 ] = 8'h9B;
ROM_MEM[556 ] = 8'h7D;
ROM_MEM[557 ] = 8'h84;
ROM_MEM[558 ] = 8'h48;
ROM_MEM[559 ] = 8'h97;
ROM_MEM[560 ] = 8'h29;
ROM_MEM[561 ] = 8'h6D;
ROM_MEM[562 ] = 8'hAA;
ROM_MEM[563 ] = 8'hA6;
ROM_MEM[564 ] = 8'h16;
ROM_MEM[565 ] = 8'h6D;
ROM_MEM[566 ] = 8'h35;
ROM_MEM[567 ] = 8'h34;
ROM_MEM[568 ] = 8'h31;
ROM_MEM[569 ] = 8'hBA;
ROM_MEM[570 ] = 8'h69;
ROM_MEM[571 ] = 8'h76;
ROM_MEM[572 ] = 8'h94;
ROM_MEM[573 ] = 8'h07;
ROM_MEM[574 ] = 8'h2A;
ROM_MEM[575 ] = 8'hEA;
ROM_MEM[576 ] = 8'hC6;
ROM_MEM[577 ] = 8'hAB;
ROM_MEM[578 ] = 8'hAB;
ROM_MEM[579 ] = 8'h41;
ROM_MEM[580 ] = 8'h37;
ROM_MEM[581 ] = 8'hCA;
ROM_MEM[582 ] = 8'hE2;
ROM_MEM[583 ] = 8'h9C;
ROM_MEM[584 ] = 8'hBA;
ROM_MEM[585 ] = 8'h04;
ROM_MEM[586 ] = 8'h5B;
ROM_MEM[587 ] = 8'h2F;
ROM_MEM[588 ] = 8'hAD;
ROM_MEM[589 ] = 8'h7D;
ROM_MEM[590 ] = 8'h8A;
ROM_MEM[591 ] = 8'h12;
ROM_MEM[592 ] = 8'h6D;
ROM_MEM[593 ] = 8'h3D;
ROM_MEM[594 ] = 8'hD3;
ROM_MEM[595 ] = 8'hF1;
ROM_MEM[596 ] = 8'hC9;
ROM_MEM[597 ] = 8'h5A;
ROM_MEM[598 ] = 8'hD4;
ROM_MEM[599 ] = 8'hD5;
ROM_MEM[600 ] = 8'hF2;
ROM_MEM[601 ] = 8'h44;
ROM_MEM[602 ] = 8'h27;
ROM_MEM[603 ] = 8'hEB;
ROM_MEM[604 ] = 8'h55;
ROM_MEM[605 ] = 8'h87;
ROM_MEM[606 ] = 8'h43;
ROM_MEM[607 ] = 8'h6B;
ROM_MEM[608 ] = 8'hAF;
ROM_MEM[609 ] = 8'hBC;
ROM_MEM[610 ] = 8'h15;
ROM_MEM[611 ] = 8'h29;
ROM_MEM[612 ] = 8'h0E;
ROM_MEM[613 ] = 8'h49;
ROM_MEM[614 ] = 8'h5C;
ROM_MEM[615 ] = 8'h8A;
ROM_MEM[616 ] = 8'h1A;
ROM_MEM[617 ] = 8'hD1;
ROM_MEM[618 ] = 8'hB4;
ROM_MEM[619 ] = 8'hD4;
ROM_MEM[620 ] = 8'hF1;
ROM_MEM[621 ] = 8'hC8;
ROM_MEM[622 ] = 8'hAB;
ROM_MEM[623 ] = 8'hE3;
ROM_MEM[624 ] = 8'hD6;
ROM_MEM[625 ] = 8'h64;
ROM_MEM[626 ] = 8'h39;
ROM_MEM[627 ] = 8'hAB;
ROM_MEM[628 ] = 8'hAE;
ROM_MEM[629 ] = 8'h4E;
ROM_MEM[630 ] = 8'hD7;
ROM_MEM[631 ] = 8'h93;
ROM_MEM[632 ] = 8'h6C;
ROM_MEM[633 ] = 8'hAF;
ROM_MEM[634 ] = 8'hBA;
ROM_MEM[635 ] = 8'h38;
ROM_MEM[636 ] = 8'h5B;
ROM_MEM[637 ] = 8'h2F;
ROM_MEM[638 ] = 8'h8E;
ROM_MEM[639 ] = 8'hB3;
ROM_MEM[640 ] = 8'h9A;
ROM_MEM[641 ] = 8'hEA;
ROM_MEM[642 ] = 8'h74;
ROM_MEM[643 ] = 8'hBD;
ROM_MEM[644 ] = 8'h28;
ROM_MEM[645 ] = 8'hCA;
ROM_MEM[646 ] = 8'h6A;
ROM_MEM[647 ] = 8'hAB;
ROM_MEM[648 ] = 8'hD3;
ROM_MEM[649 ] = 8'hB1;
ROM_MEM[650 ] = 8'hE4;
ROM_MEM[651 ] = 8'h28;
ROM_MEM[652 ] = 8'hA9;
ROM_MEM[653 ] = 8'h2D;
ROM_MEM[654 ] = 8'h8E;
ROM_MEM[655 ] = 8'h52;
ROM_MEM[656 ] = 8'hC3;
ROM_MEM[657 ] = 8'hE5;
ROM_MEM[658 ] = 8'hA6;
ROM_MEM[659 ] = 8'h26;
ROM_MEM[660 ] = 8'h2B;
ROM_MEM[661 ] = 8'hCC;
ROM_MEM[662 ] = 8'hF4;
ROM_MEM[663 ] = 8'hB4;
ROM_MEM[664 ] = 8'h13;
ROM_MEM[665 ] = 8'hDA;
ROM_MEM[666 ] = 8'hA2;
ROM_MEM[667 ] = 8'h31;
ROM_MEM[668 ] = 8'hD2;
ROM_MEM[669 ] = 8'h22;
ROM_MEM[670 ] = 8'h69;
ROM_MEM[671 ] = 8'hEB;
ROM_MEM[672 ] = 8'hAA;
ROM_MEM[673 ] = 8'hA3;
ROM_MEM[674 ] = 8'h56;
ROM_MEM[675 ] = 8'hD7;
ROM_MEM[676 ] = 8'hD6;
ROM_MEM[677 ] = 8'hA3;
ROM_MEM[678 ] = 8'hCF;
ROM_MEM[679 ] = 8'h4E;
ROM_MEM[680 ] = 8'h5A;
ROM_MEM[681 ] = 8'h22;
ROM_MEM[682 ] = 8'h9A;
ROM_MEM[683 ] = 8'h8C;
ROM_MEM[684 ] = 8'hB1;
ROM_MEM[685 ] = 8'h18;
ROM_MEM[686 ] = 8'hEA;
ROM_MEM[687 ] = 8'h30;
ROM_MEM[688 ] = 8'hCB;
ROM_MEM[689 ] = 8'h92;
ROM_MEM[690 ] = 8'hC6;
ROM_MEM[691 ] = 8'h6C;
ROM_MEM[692 ] = 8'hA8;
ROM_MEM[693 ] = 8'h02;
ROM_MEM[694 ] = 8'h7D;
ROM_MEM[695 ] = 8'h59;
ROM_MEM[696 ] = 8'h1A;
ROM_MEM[697 ] = 8'hAA;
ROM_MEM[698 ] = 8'hC3;
ROM_MEM[699 ] = 8'h70;
ROM_MEM[700 ] = 8'hB6;
ROM_MEM[701 ] = 8'hA6;
ROM_MEM[702 ] = 8'h63;
ROM_MEM[703 ] = 8'hA8;
ROM_MEM[704 ] = 8'h11;
ROM_MEM[705 ] = 8'h53;
ROM_MEM[706 ] = 8'h2B;
ROM_MEM[707 ] = 8'h56;
ROM_MEM[708 ] = 8'h8F;
ROM_MEM[709 ] = 8'hB1;
ROM_MEM[710 ] = 8'h26;
ROM_MEM[711 ] = 8'h32;
ROM_MEM[712 ] = 8'h99;
ROM_MEM[713 ] = 8'h5C;
ROM_MEM[714 ] = 8'hDD;
ROM_MEM[715 ] = 8'hA6;
ROM_MEM[716 ] = 8'h56;
ROM_MEM[717 ] = 8'hD9;
ROM_MEM[718 ] = 8'hB0;
ROM_MEM[719 ] = 8'hE2;
ROM_MEM[720 ] = 8'h75;
ROM_MEM[721 ] = 8'h59;
ROM_MEM[722 ] = 8'h6A;
ROM_MEM[723 ] = 8'h20;
ROM_MEM[724 ] = 8'h93;
ROM_MEM[725 ] = 8'hC9;
ROM_MEM[726 ] = 8'hD5;
ROM_MEM[727 ] = 8'h69;
ROM_MEM[728 ] = 8'h6B;
ROM_MEM[729 ] = 8'h59;
ROM_MEM[730 ] = 8'h54;
ROM_MEM[731 ] = 8'h59;
ROM_MEM[732 ] = 8'h52;
ROM_MEM[733 ] = 8'hB7;
ROM_MEM[734 ] = 8'hBD;
ROM_MEM[735 ] = 8'h46;
ROM_MEM[736 ] = 8'h72;
ROM_MEM[737 ] = 8'hA9;
ROM_MEM[738 ] = 8'hD8;
ROM_MEM[739 ] = 8'hD2;
ROM_MEM[740 ] = 8'h8E;
ROM_MEM[741 ] = 8'h56;
ROM_MEM[742 ] = 8'hC9;
ROM_MEM[743 ] = 8'hA5;
ROM_MEM[744 ] = 8'hAC;
ROM_MEM[745 ] = 8'hAD;
ROM_MEM[746 ] = 8'h01;
ROM_MEM[747 ] = 8'hBC;
ROM_MEM[748 ] = 8'hA5;
ROM_MEM[749 ] = 8'h56;
ROM_MEM[750 ] = 8'h40;
ROM_MEM[751 ] = 8'hB0;
ROM_MEM[752 ] = 8'h58;
ROM_MEM[753 ] = 8'h0A;
ROM_MEM[754 ] = 8'h70;
ROM_MEM[755 ] = 8'h8E;
ROM_MEM[756 ] = 8'h8A;
ROM_MEM[757 ] = 8'h01;
ROM_MEM[758 ] = 8'hDC;
ROM_MEM[759 ] = 8'h90;
ROM_MEM[760 ] = 8'h3D;
ROM_MEM[761 ] = 8'h5D;
ROM_MEM[762 ] = 8'h2D;
ROM_MEM[763 ] = 8'h4F;
ROM_MEM[764 ] = 8'h04;
ROM_MEM[765 ] = 8'h00;
ROM_MEM[766 ] = 8'hD2;
ROM_MEM[767 ] = 8'h8C;
ROM_MEM[768 ] = 8'h00;
ROM_MEM[769 ] = 8'h40;
ROM_MEM[770 ] = 8'h84;
ROM_MEM[771 ] = 8'h11;
ROM_MEM[772 ] = 8'h00;
ROM_MEM[773 ] = 8'h58;
ROM_MEM[774 ] = 8'h67;
ROM_MEM[775 ] = 8'h01;
ROM_MEM[776 ] = 8'h08;
ROM_MEM[777 ] = 8'hED;
ROM_MEM[778 ] = 8'hA6;
ROM_MEM[779 ] = 8'h00;
ROM_MEM[780 ] = 8'hE9;
ROM_MEM[781 ] = 8'hBD;
ROM_MEM[782 ] = 8'h04;
ROM_MEM[783 ] = 8'h60;
ROM_MEM[784 ] = 8'h15;
ROM_MEM[785 ] = 8'hBB;
ROM_MEM[786 ] = 8'h02;
ROM_MEM[787 ] = 8'hBC;
ROM_MEM[788 ] = 8'h64;
ROM_MEM[789 ] = 8'h17;
ROM_MEM[790 ] = 8'h80;
ROM_MEM[791 ] = 8'h36;
ROM_MEM[792 ] = 8'hA2;
ROM_MEM[793 ] = 8'h02;
ROM_MEM[794 ] = 8'hD0;
ROM_MEM[795 ] = 8'h5A;
ROM_MEM[796 ] = 8'h35;
ROM_MEM[797 ] = 8'h35;
ROM_MEM[798 ] = 8'h59;
ROM_MEM[799 ] = 8'h6A;
ROM_MEM[800 ] = 8'hB1;
ROM_MEM[801 ] = 8'h47;
ROM_MEM[802 ] = 8'hEA;
ROM_MEM[803 ] = 8'hD2;
ROM_MEM[804 ] = 8'h79;
ROM_MEM[805 ] = 8'h19;
ROM_MEM[806 ] = 8'h2B;
ROM_MEM[807 ] = 8'h69;
ROM_MEM[808 ] = 8'h8E;
ROM_MEM[809 ] = 8'h5A;
ROM_MEM[810 ] = 8'h6B;
ROM_MEM[811 ] = 8'h4D;
ROM_MEM[812 ] = 8'hAE;
ROM_MEM[813 ] = 8'h54;
ROM_MEM[814 ] = 8'hB8;
ROM_MEM[815 ] = 8'h6A;
ROM_MEM[816 ] = 8'hAD;
ROM_MEM[817 ] = 8'h71;
ROM_MEM[818 ] = 8'hB9;
ROM_MEM[819 ] = 8'h56;
ROM_MEM[820 ] = 8'hEA;
ROM_MEM[821 ] = 8'hAA;
ROM_MEM[822 ] = 8'h75;
ROM_MEM[823 ] = 8'hC1;
ROM_MEM[824 ] = 8'hDB;
ROM_MEM[825 ] = 8'hB0;
ROM_MEM[826 ] = 8'hF1;
ROM_MEM[827 ] = 8'hA6;
ROM_MEM[828 ] = 8'hD6;
ROM_MEM[829 ] = 8'hA5;
ROM_MEM[830 ] = 8'h1A;
ROM_MEM[831 ] = 8'h43;
ROM_MEM[832 ] = 8'h64;
ROM_MEM[833 ] = 8'h89;
ROM_MEM[834 ] = 8'h7B;
ROM_MEM[835 ] = 8'h67;
ROM_MEM[836 ] = 8'h80;
ROM_MEM[837 ] = 8'h0C;
ROM_MEM[838 ] = 8'hC5;
ROM_MEM[839 ] = 8'h0C;
ROM_MEM[840 ] = 8'h50;
ROM_MEM[841 ] = 8'h20;
ROM_MEM[842 ] = 8'h73;
ROM_MEM[843 ] = 8'h19;
ROM_MEM[844 ] = 8'h8B;
ROM_MEM[845 ] = 8'h34;
ROM_MEM[846 ] = 8'h49;
ROM_MEM[847 ] = 8'hF5;
ROM_MEM[848 ] = 8'hB4;
ROM_MEM[849 ] = 8'h6D;
ROM_MEM[850 ] = 8'hCE;
ROM_MEM[851 ] = 8'h5A;
ROM_MEM[852 ] = 8'hDC;
ROM_MEM[853 ] = 8'hC5;
ROM_MEM[854 ] = 8'h5B;
ROM_MEM[855 ] = 8'h8F;
ROM_MEM[856 ] = 8'h75;
ROM_MEM[857 ] = 8'hC7;
ROM_MEM[858 ] = 8'h54;
ROM_MEM[859 ] = 8'h53;
ROM_MEM[860 ] = 8'h95;
ROM_MEM[861 ] = 8'hEA;
ROM_MEM[862 ] = 8'h80;
ROM_MEM[863 ] = 8'h21;
ROM_MEM[864 ] = 8'h81;
ROM_MEM[865 ] = 8'h13;
ROM_MEM[866 ] = 8'h30;
ROM_MEM[867 ] = 8'h25;
ROM_MEM[868 ] = 8'h51;
ROM_MEM[869 ] = 8'h02;
ROM_MEM[870 ] = 8'hA6;
ROM_MEM[871 ] = 8'h43;
ROM_MEM[872 ] = 8'h29;
ROM_MEM[873 ] = 8'hC0;
ROM_MEM[874 ] = 8'h8C;
ROM_MEM[875 ] = 8'h2C;
ROM_MEM[876 ] = 8'h05;
ROM_MEM[877 ] = 8'h98;
ROM_MEM[878 ] = 8'h41;
ROM_MEM[879 ] = 8'h29;
ROM_MEM[880 ] = 8'h01;
ROM_MEM[881 ] = 8'hCB;
ROM_MEM[882 ] = 8'h12;
ROM_MEM[883 ] = 8'h2A;
ROM_MEM[884 ] = 8'h20;
ROM_MEM[885 ] = 8'h50;
ROM_MEM[886 ] = 8'h32;
ROM_MEM[887 ] = 8'h02;
ROM_MEM[888 ] = 8'h48;
ROM_MEM[889 ] = 8'h8C;
ROM_MEM[890 ] = 8'h49;
ROM_MEM[891 ] = 8'h00;
ROM_MEM[892 ] = 8'h40;
ROM_MEM[893 ] = 8'hC5;
ROM_MEM[894 ] = 8'h0C;
ROM_MEM[895 ] = 8'h50;
ROM_MEM[896 ] = 8'h02;
ROM_MEM[897 ] = 8'h78;
ROM_MEM[898 ] = 8'h00;
ROM_MEM[899 ] = 8'h5A;
ROM_MEM[900 ] = 8'h60;
ROM_MEM[901 ] = 8'h1C;
ROM_MEM[902 ] = 8'hB1;
ROM_MEM[903 ] = 8'hCF;
ROM_MEM[904 ] = 8'h1E;
ROM_MEM[905 ] = 8'hAA;
ROM_MEM[906 ] = 8'h9E;
ROM_MEM[907 ] = 8'h74;
ROM_MEM[908 ] = 8'h44;
ROM_MEM[909 ] = 8'h66;
ROM_MEM[910 ] = 8'h5A;
ROM_MEM[911 ] = 8'h48;
ROM_MEM[912 ] = 8'hA4;
ROM_MEM[913 ] = 8'hBB;
ROM_MEM[914 ] = 8'h95;
ROM_MEM[915 ] = 8'h44;
ROM_MEM[916 ] = 8'hAB;
ROM_MEM[917 ] = 8'h2B;
ROM_MEM[918 ] = 8'hC1;
ROM_MEM[919 ] = 8'h69;
ROM_MEM[920 ] = 8'h4F;
ROM_MEM[921 ] = 8'h9E;
ROM_MEM[922 ] = 8'h8C;
ROM_MEM[923 ] = 8'hAD;
ROM_MEM[924 ] = 8'h3A;
ROM_MEM[925 ] = 8'h75;
ROM_MEM[926 ] = 8'h3E;
ROM_MEM[927 ] = 8'h6D;
ROM_MEM[928 ] = 8'h51;
ROM_MEM[929 ] = 8'hBA;
ROM_MEM[930 ] = 8'h5E;
ROM_MEM[931 ] = 8'h98;
ROM_MEM[932 ] = 8'hE7;
ROM_MEM[933 ] = 8'hAC;
ROM_MEM[934 ] = 8'h55;
ROM_MEM[935 ] = 8'hEB;
ROM_MEM[936 ] = 8'hC6;
ROM_MEM[937 ] = 8'h40;
ROM_MEM[938 ] = 8'hD2;
ROM_MEM[939 ] = 8'hB5;
ROM_MEM[940 ] = 8'h15;
ROM_MEM[941 ] = 8'h6D;
ROM_MEM[942 ] = 8'hEB;
ROM_MEM[943 ] = 8'h05;
ROM_MEM[944 ] = 8'h49;
ROM_MEM[945 ] = 8'hC6;
ROM_MEM[946 ] = 8'h5E;
ROM_MEM[947 ] = 8'h95;
ROM_MEM[948 ] = 8'hAD;
ROM_MEM[949 ] = 8'h35;
ROM_MEM[950 ] = 8'hC9;
ROM_MEM[951 ] = 8'h2E;
ROM_MEM[952 ] = 8'h5B;
ROM_MEM[953 ] = 8'h32;
ROM_MEM[954 ] = 8'h3E;
ROM_MEM[955 ] = 8'hC6;
ROM_MEM[956 ] = 8'hA4;
ROM_MEM[957 ] = 8'h24;
ROM_MEM[958 ] = 8'hED;
ROM_MEM[959 ] = 8'h45;
ROM_MEM[960 ] = 8'h63;
ROM_MEM[961 ] = 8'h46;
ROM_MEM[962 ] = 8'hB8;
ROM_MEM[963 ] = 8'hE4;
ROM_MEM[964 ] = 8'hB4;
ROM_MEM[965 ] = 8'h17;
ROM_MEM[966 ] = 8'h8D;
ROM_MEM[967 ] = 8'h91;
ROM_MEM[968 ] = 8'h15;
ROM_MEM[969 ] = 8'h92;
ROM_MEM[970 ] = 8'hC3;
ROM_MEM[971 ] = 8'h5E;
ROM_MEM[972 ] = 8'h35;
ROM_MEM[973 ] = 8'h78;
ROM_MEM[974 ] = 8'h65;
ROM_MEM[975 ] = 8'h99;
ROM_MEM[976 ] = 8'h76;
ROM_MEM[977 ] = 8'h7B;
ROM_MEM[978 ] = 8'hE6;
ROM_MEM[979 ] = 8'h1C;
ROM_MEM[980 ] = 8'h93;
ROM_MEM[981 ] = 8'h2E;
ROM_MEM[982 ] = 8'h51;
ROM_MEM[983 ] = 8'h00;
ROM_MEM[984 ] = 8'hCC;
ROM_MEM[985 ] = 8'h45;
ROM_MEM[986 ] = 8'h2A;
ROM_MEM[987 ] = 8'h40;
ROM_MEM[988 ] = 8'h73;
ROM_MEM[989 ] = 8'h2D;
ROM_MEM[990 ] = 8'h03;
ROM_MEM[991 ] = 8'h04;
ROM_MEM[992 ] = 8'hC5;
ROM_MEM[993 ] = 8'h1D;
ROM_MEM[994 ] = 8'hFA;
ROM_MEM[995 ] = 8'hEE;
ROM_MEM[996 ] = 8'h59;
ROM_MEM[997 ] = 8'h55;
ROM_MEM[998 ] = 8'h35;
ROM_MEM[999 ] = 8'h0D;
ROM_MEM[1000] = 8'h03;
ROM_MEM[1001] = 8'hB0;
ROM_MEM[1002] = 8'h94;
ROM_MEM[1003] = 8'h6E;
ROM_MEM[1004] = 8'h7B;
ROM_MEM[1005] = 8'h73;
ROM_MEM[1006] = 8'hE4;
ROM_MEM[1007] = 8'hE6;
ROM_MEM[1008] = 8'hDE;
ROM_MEM[1009] = 8'hB6;
ROM_MEM[1010] = 8'hED;
ROM_MEM[1011] = 8'hD5;
ROM_MEM[1012] = 8'hA2;
ROM_MEM[1013] = 8'h7B;
ROM_MEM[1014] = 8'h7B;
ROM_MEM[1015] = 8'hDB;
ROM_MEM[1016] = 8'hB2;
ROM_MEM[1017] = 8'h67;
ROM_MEM[1018] = 8'hC9;
ROM_MEM[1019] = 8'h35;
ROM_MEM[1020] = 8'hE5;
ROM_MEM[1021] = 8'h49;
ROM_MEM[1022] = 8'h04;
ROM_MEM[1023] = 8'h60;
ROM_MEM[1024] = 8'hA0;
ROM_MEM[1025] = 8'h86;
ROM_MEM[1026] = 8'h00;
ROM_MEM[1027] = 8'h3C;
ROM_MEM[1028] = 8'h64;
ROM_MEM[1029] = 8'h31;
ROM_MEM[1030] = 8'h40;
ROM_MEM[1031] = 8'h17;
ROM_MEM[1032] = 8'hA0;
ROM_MEM[1033] = 8'h02;
ROM_MEM[1034] = 8'hE0;
ROM_MEM[1035] = 8'hDE;
ROM_MEM[1036] = 8'hD4;
ROM_MEM[1037] = 8'h95;
ROM_MEM[1038] = 8'h5E;
ROM_MEM[1039] = 8'h45;
ROM_MEM[1040] = 8'h99;
ROM_MEM[1041] = 8'h68;
ROM_MEM[1042] = 8'hDA;
ROM_MEM[1043] = 8'h94;
ROM_MEM[1044] = 8'h27;
ROM_MEM[1045] = 8'h2D;
ROM_MEM[1046] = 8'hE5;
ROM_MEM[1047] = 8'hAA;
ROM_MEM[1048] = 8'h8D;
ROM_MEM[1049] = 8'h53;
ROM_MEM[1050] = 8'h55;
ROM_MEM[1051] = 8'h0C;
ROM_MEM[1052] = 8'hBA;
ROM_MEM[1053] = 8'hAB;
ROM_MEM[1054] = 8'hC9;
ROM_MEM[1055] = 8'h4D;
ROM_MEM[1056] = 8'h4D;
ROM_MEM[1057] = 8'h31;
ROM_MEM[1058] = 8'hE8;
ROM_MEM[1059] = 8'hEC;
ROM_MEM[1060] = 8'hE1;
ROM_MEM[1061] = 8'hCE;
ROM_MEM[1062] = 8'h0D;
ROM_MEM[1063] = 8'h45;
ROM_MEM[1064] = 8'hB0;
ROM_MEM[1065] = 8'hB8;
ROM_MEM[1066] = 8'h55;
ROM_MEM[1067] = 8'h12;
ROM_MEM[1068] = 8'hB3;
ROM_MEM[1069] = 8'h55;
ROM_MEM[1070] = 8'hCE;
ROM_MEM[1071] = 8'hA2;
ROM_MEM[1072] = 8'h9E;
ROM_MEM[1073] = 8'h49;
ROM_MEM[1074] = 8'h1E;
ROM_MEM[1075] = 8'h00;
ROM_MEM[1076] = 8'h44;
ROM_MEM[1077] = 8'h15;
ROM_MEM[1078] = 8'h21;
ROM_MEM[1079] = 8'hD4;
ROM_MEM[1080] = 8'h21;
ROM_MEM[1081] = 8'h2D;
ROM_MEM[1082] = 8'h2B;
ROM_MEM[1083] = 8'h15;
ROM_MEM[1084] = 8'h0F;
ROM_MEM[1085] = 8'h5F;
ROM_MEM[1086] = 8'h17;
ROM_MEM[1087] = 8'h8F;
ROM_MEM[1088] = 8'hAE;
ROM_MEM[1089] = 8'hB4;
ROM_MEM[1090] = 8'hB5;
ROM_MEM[1091] = 8'h3C;
ROM_MEM[1092] = 8'hD3;
ROM_MEM[1093] = 8'h22;
ROM_MEM[1094] = 8'h37;
ROM_MEM[1095] = 8'h32;
ROM_MEM[1096] = 8'hF2;
ROM_MEM[1097] = 8'h71;
ROM_MEM[1098] = 8'h7D;
ROM_MEM[1099] = 8'hB2;
ROM_MEM[1100] = 8'hDC;
ROM_MEM[1101] = 8'h6C;
ROM_MEM[1102] = 8'h2B;
ROM_MEM[1103] = 8'hC7;
ROM_MEM[1104] = 8'h4D;
ROM_MEM[1105] = 8'hD6;
ROM_MEM[1106] = 8'hA2;
ROM_MEM[1107] = 8'h72;
ROM_MEM[1108] = 8'hAD;
ROM_MEM[1109] = 8'h14;
ROM_MEM[1110] = 8'h3F;
ROM_MEM[1111] = 8'h5A;
ROM_MEM[1112] = 8'hF1;
ROM_MEM[1113] = 8'hCC;
ROM_MEM[1114] = 8'hA6;
ROM_MEM[1115] = 8'h54;
ROM_MEM[1116] = 8'hC2;
ROM_MEM[1117] = 8'h60;
ROM_MEM[1118] = 8'h54;
ROM_MEM[1119] = 8'hD3;
ROM_MEM[1120] = 8'h42;
ROM_MEM[1121] = 8'h4A;
ROM_MEM[1122] = 8'h88;
ROM_MEM[1123] = 8'h32;
ROM_MEM[1124] = 8'h75;
ROM_MEM[1125] = 8'h35;
ROM_MEM[1126] = 8'h4F;
ROM_MEM[1127] = 8'hD3;
ROM_MEM[1128] = 8'h0C;
ROM_MEM[1129] = 8'hA0;
ROM_MEM[1130] = 8'h3A;
ROM_MEM[1131] = 8'h8C;
ROM_MEM[1132] = 8'h01;
ROM_MEM[1133] = 8'h4C;
ROM_MEM[1134] = 8'h6A;
ROM_MEM[1135] = 8'h08;
ROM_MEM[1136] = 8'h80;
ROM_MEM[1137] = 8'h4B;
ROM_MEM[1138] = 8'h37;
ROM_MEM[1139] = 8'h01;
ROM_MEM[1140] = 8'h28;
ROM_MEM[1141] = 8'hA6;
ROM_MEM[1142] = 8'hB2;
ROM_MEM[1143] = 8'h74;
ROM_MEM[1144] = 8'h3F;
ROM_MEM[1145] = 8'hCD;
ROM_MEM[1146] = 8'h43;
ROM_MEM[1147] = 8'h3A;
ROM_MEM[1148] = 8'hEC;
ROM_MEM[1149] = 8'h30;
ROM_MEM[1150] = 8'hFC;
ROM_MEM[1151] = 8'h51;
ROM_MEM[1152] = 8'h8F;
ROM_MEM[1153] = 8'hE8;
ROM_MEM[1154] = 8'h4A;
ROM_MEM[1155] = 8'hCB;
ROM_MEM[1156] = 8'h0C;
ROM_MEM[1157] = 8'hDB;
ROM_MEM[1158] = 8'hDC;
ROM_MEM[1159] = 8'h7D;
ROM_MEM[1160] = 8'hAA;
ROM_MEM[1161] = 8'h2E;
ROM_MEM[1162] = 8'h33;
ROM_MEM[1163] = 8'h6C;
ROM_MEM[1164] = 8'h89;
ROM_MEM[1165] = 8'h88;
ROM_MEM[1166] = 8'h09;
ROM_MEM[1167] = 8'hBB;
ROM_MEM[1168] = 8'hAC;
ROM_MEM[1169] = 8'hB0;
ROM_MEM[1170] = 8'hC5;
ROM_MEM[1171] = 8'h33;
ROM_MEM[1172] = 8'h26;
ROM_MEM[1173] = 8'hEC;
ROM_MEM[1174] = 8'hB2;
ROM_MEM[1175] = 8'hC2;
ROM_MEM[1176] = 8'hB6;
ROM_MEM[1177] = 8'hF0;
ROM_MEM[1178] = 8'h68;
ROM_MEM[1179] = 8'hB3;
ROM_MEM[1180] = 8'hCB;
ROM_MEM[1181] = 8'h0E;
ROM_MEM[1182] = 8'hCB;
ROM_MEM[1183] = 8'h22;
ROM_MEM[1184] = 8'hBC;
ROM_MEM[1185] = 8'hCD;
ROM_MEM[1186] = 8'h2D;
ROM_MEM[1187] = 8'h3B;
ROM_MEM[1188] = 8'h76;
ROM_MEM[1189] = 8'h2D;
ROM_MEM[1190] = 8'hCB;
ROM_MEM[1191] = 8'h96;
ROM_MEM[1192] = 8'h7A;
ROM_MEM[1193] = 8'hDC;
ROM_MEM[1194] = 8'h54;
ROM_MEM[1195] = 8'hB8;
ROM_MEM[1196] = 8'hAC;
ROM_MEM[1197] = 8'h4B;
ROM_MEM[1198] = 8'hCE;
ROM_MEM[1199] = 8'hF2;
ROM_MEM[1200] = 8'h82;
ROM_MEM[1201] = 8'hD7;
ROM_MEM[1202] = 8'h29;
ROM_MEM[1203] = 8'h6F;
ROM_MEM[1204] = 8'hB9;
ROM_MEM[1205] = 8'h25;
ROM_MEM[1206] = 8'h0C;
ROM_MEM[1207] = 8'h4E;
ROM_MEM[1208] = 8'h3C;
ROM_MEM[1209] = 8'hBD;
ROM_MEM[1210] = 8'h22;
ROM_MEM[1211] = 8'hA5;
ROM_MEM[1212] = 8'h28;
ROM_MEM[1213] = 8'h29;
ROM_MEM[1214] = 8'h37;
ROM_MEM[1215] = 8'h55;
ROM_MEM[1216] = 8'hB3;
ROM_MEM[1217] = 8'h62;
ROM_MEM[1218] = 8'h00;
ROM_MEM[1219] = 8'hA7;
ROM_MEM[1220] = 8'h42;
ROM_MEM[1221] = 8'h15;
ROM_MEM[1222] = 8'hA0;
ROM_MEM[1223] = 8'h48;
ROM_MEM[1224] = 8'h39;
ROM_MEM[1225] = 8'h01;
ROM_MEM[1226] = 8'h80;
ROM_MEM[1227] = 8'h37;
ROM_MEM[1228] = 8'h53;
ROM_MEM[1229] = 8'h80;
ROM_MEM[1230] = 8'h15;
ROM_MEM[1231] = 8'h69;
ROM_MEM[1232] = 8'hCB;
ROM_MEM[1233] = 8'h4F;
ROM_MEM[1234] = 8'hDA;
ROM_MEM[1235] = 8'h74;
ROM_MEM[1236] = 8'h33;
ROM_MEM[1237] = 8'h8D;
ROM_MEM[1238] = 8'hAC;
ROM_MEM[1239] = 8'h20;
ROM_MEM[1240] = 8'h5B;
ROM_MEM[1241] = 8'hF6;
ROM_MEM[1242] = 8'hAD;
ROM_MEM[1243] = 8'h36;
ROM_MEM[1244] = 8'hB2;
ROM_MEM[1245] = 8'hC2;
ROM_MEM[1246] = 8'h62;
ROM_MEM[1247] = 8'h39;
ROM_MEM[1248] = 8'h2A;
ROM_MEM[1249] = 8'h87;
ROM_MEM[1250] = 8'hF2;
ROM_MEM[1251] = 8'h89;
ROM_MEM[1252] = 8'hAA;
ROM_MEM[1253] = 8'h67;
ROM_MEM[1254] = 8'hAB;
ROM_MEM[1255] = 8'h5C;
ROM_MEM[1256] = 8'h29;
ROM_MEM[1257] = 8'h27;
ROM_MEM[1258] = 8'hAA;
ROM_MEM[1259] = 8'h51;
ROM_MEM[1260] = 8'hCC;
ROM_MEM[1261] = 8'h6B;
ROM_MEM[1262] = 8'hA9;
ROM_MEM[1263] = 8'hAC;
ROM_MEM[1264] = 8'hB8;
ROM_MEM[1265] = 8'h44;
ROM_MEM[1266] = 8'h51;
ROM_MEM[1267] = 8'hEF;
ROM_MEM[1268] = 8'h95;
ROM_MEM[1269] = 8'h52;
ROM_MEM[1270] = 8'h12;
ROM_MEM[1271] = 8'hE5;
ROM_MEM[1272] = 8'h32;
ROM_MEM[1273] = 8'h4A;
ROM_MEM[1274] = 8'hC2;
ROM_MEM[1275] = 8'hCA;
ROM_MEM[1276] = 8'h4A;
ROM_MEM[1277] = 8'hB2;
ROM_MEM[1278] = 8'h14;
ROM_MEM[1279] = 8'hAF;
ROM_MEM[1280] = 8'h1C;
ROM_MEM[1281] = 8'h29;
ROM_MEM[1282] = 8'h2B;
ROM_MEM[1283] = 8'hA9;
ROM_MEM[1284] = 8'h86;
ROM_MEM[1285] = 8'hA2;
ROM_MEM[1286] = 8'h22;
ROM_MEM[1287] = 8'h94;
ROM_MEM[1288] = 8'h8C;
ROM_MEM[1289] = 8'h24;
ROM_MEM[1290] = 8'h2B;
ROM_MEM[1291] = 8'hCA;
ROM_MEM[1292] = 8'hD3;
ROM_MEM[1293] = 8'h90;
ROM_MEM[1294] = 8'h5A;
ROM_MEM[1295] = 8'h52;
ROM_MEM[1296] = 8'h65;
ROM_MEM[1297] = 8'hCB;
ROM_MEM[1298] = 8'h8B;
ROM_MEM[1299] = 8'hDD;
ROM_MEM[1300] = 8'h76;
ROM_MEM[1301] = 8'hC8;
ROM_MEM[1302] = 8'h84;
ROM_MEM[1303] = 8'hA9;
ROM_MEM[1304] = 8'h68;
ROM_MEM[1305] = 8'h33;
ROM_MEM[1306] = 8'hC7;
ROM_MEM[1307] = 8'h21;
ROM_MEM[1308] = 8'hF7;
ROM_MEM[1309] = 8'hDA;
ROM_MEM[1310] = 8'h3D;
ROM_MEM[1311] = 8'hDD;
ROM_MEM[1312] = 8'hE2;
ROM_MEM[1313] = 8'h8C;
ROM_MEM[1314] = 8'hCC;
ROM_MEM[1315] = 8'h77;
ROM_MEM[1316] = 8'h0B;
ROM_MEM[1317] = 8'h8F;
ROM_MEM[1318] = 8'h29;
ROM_MEM[1319] = 8'h3C;
ROM_MEM[1320] = 8'h52;
ROM_MEM[1321] = 8'hDF;
ROM_MEM[1322] = 8'hB5;
ROM_MEM[1323] = 8'h34;
ROM_MEM[1324] = 8'h37;
ROM_MEM[1325] = 8'hCC;
ROM_MEM[1326] = 8'h48;
ROM_MEM[1327] = 8'hC3;
ROM_MEM[1328] = 8'hD4;
ROM_MEM[1329] = 8'h92;
ROM_MEM[1330] = 8'h5E;
ROM_MEM[1331] = 8'hCB;
ROM_MEM[1332] = 8'h2D;
ROM_MEM[1333] = 8'h09;
ROM_MEM[1334] = 8'h5B;
ROM_MEM[1335] = 8'hCA;
ROM_MEM[1336] = 8'hA6;
ROM_MEM[1337] = 8'hAD;
ROM_MEM[1338] = 8'h8C;
ROM_MEM[1339] = 8'h24;
ROM_MEM[1340] = 8'h2C;
ROM_MEM[1341] = 8'h4D;
ROM_MEM[1342] = 8'hAB;
ROM_MEM[1343] = 8'hB1;
ROM_MEM[1344] = 8'h32;
ROM_MEM[1345] = 8'hE2;
ROM_MEM[1346] = 8'h30;
ROM_MEM[1347] = 8'hAC;
ROM_MEM[1348] = 8'hA4;
ROM_MEM[1349] = 8'hDB;
ROM_MEM[1350] = 8'hCA;
ROM_MEM[1351] = 8'h8A;
ROM_MEM[1352] = 8'h43;
ROM_MEM[1353] = 8'hF5;
ROM_MEM[1354] = 8'hE1;
ROM_MEM[1355] = 8'h2E;
ROM_MEM[1356] = 8'h3B;
ROM_MEM[1357] = 8'h27;
ROM_MEM[1358] = 8'h8E;
ROM_MEM[1359] = 8'hC5;
ROM_MEM[1360] = 8'hDA;
ROM_MEM[1361] = 8'hB2;
ROM_MEM[1362] = 8'h65;
ROM_MEM[1363] = 8'hAF;
ROM_MEM[1364] = 8'h38;
ROM_MEM[1365] = 8'h06;
ROM_MEM[1366] = 8'h19;
ROM_MEM[1367] = 8'hAF;
ROM_MEM[1368] = 8'h96;
ROM_MEM[1369] = 8'hBC;
ROM_MEM[1370] = 8'hE2;
ROM_MEM[1371] = 8'hE8;
ROM_MEM[1372] = 8'h64;
ROM_MEM[1373] = 8'h7D;
ROM_MEM[1374] = 8'h92;
ROM_MEM[1375] = 8'h4E;
ROM_MEM[1376] = 8'h8B;
ROM_MEM[1377] = 8'hB3;
ROM_MEM[1378] = 8'hC7;
ROM_MEM[1379] = 8'h8A;
ROM_MEM[1380] = 8'h6A;
ROM_MEM[1381] = 8'hB1;
ROM_MEM[1382] = 8'h2E;
ROM_MEM[1383] = 8'h0E;
ROM_MEM[1384] = 8'hC2;
ROM_MEM[1385] = 8'hC4;
ROM_MEM[1386] = 8'h22;
ROM_MEM[1387] = 8'h1C;
ROM_MEM[1388] = 8'hBB;
ROM_MEM[1389] = 8'hB8;
ROM_MEM[1390] = 8'h08;
ROM_MEM[1391] = 8'h37;
ROM_MEM[1392] = 8'h73;
ROM_MEM[1393] = 8'h93;
ROM_MEM[1394] = 8'hFD;
ROM_MEM[1395] = 8'h00;
ROM_MEM[1396] = 8'hF7;
ROM_MEM[1397] = 8'hA9;
ROM_MEM[1398] = 8'hBA;
ROM_MEM[1399] = 8'h04;
ROM_MEM[1400] = 8'hA0;
ROM_MEM[1401] = 8'h65;
ROM_MEM[1402] = 8'h32;
ROM_MEM[1403] = 8'hB8;
ROM_MEM[1404] = 8'h49;
ROM_MEM[1405] = 8'hB9;
ROM_MEM[1406] = 8'h45;
ROM_MEM[1407] = 8'hB6;
ROM_MEM[1408] = 8'h45;
ROM_MEM[1409] = 8'h03;
ROM_MEM[1410] = 8'h60;
ROM_MEM[1411] = 8'h99;
ROM_MEM[1412] = 8'h21;
ROM_MEM[1413] = 8'h00;
ROM_MEM[1414] = 8'h4B;
ROM_MEM[1415] = 8'h34;
ROM_MEM[1416] = 8'h14;
ROM_MEM[1417] = 8'h10;
ROM_MEM[1418] = 8'hA1;
ROM_MEM[1419] = 8'hBA;
ROM_MEM[1420] = 8'h00;
ROM_MEM[1421] = 8'h0C;
ROM_MEM[1422] = 8'hF3;
ROM_MEM[1423] = 8'h66;
ROM_MEM[1424] = 8'h00;
ROM_MEM[1425] = 8'hF1;
ROM_MEM[1426] = 8'h95;
ROM_MEM[1427] = 8'h04;
ROM_MEM[1428] = 8'h40;
ROM_MEM[1429] = 8'hA9;
ROM_MEM[1430] = 8'h23;
ROM_MEM[1431] = 8'h78;
ROM_MEM[1432] = 8'h31;
ROM_MEM[1433] = 8'hA8;
ROM_MEM[1434] = 8'h7A;
ROM_MEM[1435] = 8'hBA;
ROM_MEM[1436] = 8'h93;
ROM_MEM[1437] = 8'hE6;
ROM_MEM[1438] = 8'hC4;
ROM_MEM[1439] = 8'h8A;
ROM_MEM[1440] = 8'h95;
ROM_MEM[1441] = 8'h9A;
ROM_MEM[1442] = 8'h8D;
ROM_MEM[1443] = 8'h96;
ROM_MEM[1444] = 8'h13;
ROM_MEM[1445] = 8'h13;
ROM_MEM[1446] = 8'h77;
ROM_MEM[1447] = 8'hFB;
ROM_MEM[1448] = 8'h24;
ROM_MEM[1449] = 8'h3E;
ROM_MEM[1450] = 8'h6E;
ROM_MEM[1451] = 8'h8A;
ROM_MEM[1452] = 8'h94;
ROM_MEM[1453] = 8'h95;
ROM_MEM[1454] = 8'hE7;
ROM_MEM[1455] = 8'h28;
ROM_MEM[1456] = 8'h04;
ROM_MEM[1457] = 8'hD1;
ROM_MEM[1458] = 8'h72;
ROM_MEM[1459] = 8'h44;
ROM_MEM[1460] = 8'hA4;
ROM_MEM[1461] = 8'h48;
ROM_MEM[1462] = 8'h13;
ROM_MEM[1463] = 8'h1A;
ROM_MEM[1464] = 8'hD9;
ROM_MEM[1465] = 8'hE1;
ROM_MEM[1466] = 8'hE1;
ROM_MEM[1467] = 8'h94;
ROM_MEM[1468] = 8'h19;
ROM_MEM[1469] = 8'h00;
ROM_MEM[1470] = 8'h8D;
ROM_MEM[1471] = 8'h27;
ROM_MEM[1472] = 8'h02;
ROM_MEM[1473] = 8'h3C;
ROM_MEM[1474] = 8'h13;
ROM_MEM[1475] = 8'h41;
ROM_MEM[1476] = 8'h40;
ROM_MEM[1477] = 8'h24;
ROM_MEM[1478] = 8'hA2;
ROM_MEM[1479] = 8'h08;
ROM_MEM[1480] = 8'h48;
ROM_MEM[1481] = 8'h94;
ROM_MEM[1482] = 8'h95;
ROM_MEM[1483] = 8'h00;
ROM_MEM[1484] = 8'h95;
ROM_MEM[1485] = 8'hA9;
ROM_MEM[1486] = 8'h0C;
ROM_MEM[1487] = 8'hC7;
ROM_MEM[1488] = 8'hCF;
ROM_MEM[1489] = 8'h70;
ROM_MEM[1490] = 8'hB7;
ROM_MEM[1491] = 8'hAC;
ROM_MEM[1492] = 8'hB2;
ROM_MEM[1493] = 8'h5C;
ROM_MEM[1494] = 8'h7F;
ROM_MEM[1495] = 8'h23;
ROM_MEM[1496] = 8'h4D;
ROM_MEM[1497] = 8'hAB;
ROM_MEM[1498] = 8'hCA;
ROM_MEM[1499] = 8'hF2;
ROM_MEM[1500] = 8'hC3;
ROM_MEM[1501] = 8'hD3;
ROM_MEM[1502] = 8'hB0;
ROM_MEM[1503] = 8'h9C;
ROM_MEM[1504] = 8'h24;
ROM_MEM[1505] = 8'h2B;
ROM_MEM[1506] = 8'h0C;
ROM_MEM[1507] = 8'hD7;
ROM_MEM[1508] = 8'h4B;
ROM_MEM[1509] = 8'h62;
ROM_MEM[1510] = 8'hE2;
ROM_MEM[1511] = 8'hAC;
ROM_MEM[1512] = 8'h28;
ROM_MEM[1513] = 8'h6C;
ROM_MEM[1514] = 8'h4F;
ROM_MEM[1515] = 8'hF3;
ROM_MEM[1516] = 8'h8E;
ROM_MEM[1517] = 8'hB3;
ROM_MEM[1518] = 8'hE2;
ROM_MEM[1519] = 8'hB0;
ROM_MEM[1520] = 8'hAC;
ROM_MEM[1521] = 8'hA5;
ROM_MEM[1522] = 8'hC6;
ROM_MEM[1523] = 8'hCE;
ROM_MEM[1524] = 8'h4A;
ROM_MEM[1525] = 8'h42;
ROM_MEM[1526] = 8'hF7;
ROM_MEM[1527] = 8'h91;
ROM_MEM[1528] = 8'h6C;
ROM_MEM[1529] = 8'hDB;
ROM_MEM[1530] = 8'h2B;
ROM_MEM[1531] = 8'h8B;
ROM_MEM[1532] = 8'hD9;
ROM_MEM[1533] = 8'h46;
ROM_MEM[1534] = 8'h73;
ROM_MEM[1535] = 8'h6C;
ROM_MEM[1536] = 8'hAF;
ROM_MEM[1537] = 8'h3C;
ROM_MEM[1538] = 8'h66;
ROM_MEM[1539] = 8'h1B;
ROM_MEM[1540] = 8'hEB;
ROM_MEM[1541] = 8'hB6;
ROM_MEM[1542] = 8'hBD;
ROM_MEM[1543] = 8'h8A;
ROM_MEM[1544] = 8'h90;
ROM_MEM[1545] = 8'h74;
ROM_MEM[1546] = 8'hB4;
ROM_MEM[1547] = 8'hC7;
ROM_MEM[1548] = 8'h76;
ROM_MEM[1549] = 8'hAA;
ROM_MEM[1550] = 8'hA2;
ROM_MEM[1551] = 8'hE7;
ROM_MEM[1552] = 8'h72;
ROM_MEM[1553] = 8'hC9;
ROM_MEM[1554] = 8'h5A;
ROM_MEM[1555] = 8'h29;
ROM_MEM[1556] = 8'hF1;
ROM_MEM[1557] = 8'hD1;
ROM_MEM[1558] = 8'hCC;
ROM_MEM[1559] = 8'hDD;
ROM_MEM[1560] = 8'h63;
ROM_MEM[1561] = 8'hB5;
ROM_MEM[1562] = 8'h38;
ROM_MEM[1563] = 8'h64;
ROM_MEM[1564] = 8'hCD;
ROM_MEM[1565] = 8'hD4;
ROM_MEM[1566] = 8'h8A;
ROM_MEM[1567] = 8'h34;
ROM_MEM[1568] = 8'h62;
ROM_MEM[1569] = 8'h5F;
ROM_MEM[1570] = 8'hA5;
ROM_MEM[1571] = 8'h2D;
ROM_MEM[1572] = 8'hC6;
ROM_MEM[1573] = 8'h4A;
ROM_MEM[1574] = 8'h4B;
ROM_MEM[1575] = 8'hBC;
ROM_MEM[1576] = 8'hB5;
ROM_MEM[1577] = 8'h48;
ROM_MEM[1578] = 8'hF6;
ROM_MEM[1579] = 8'hC6;
ROM_MEM[1580] = 8'h25;
ROM_MEM[1581] = 8'hB2;
ROM_MEM[1582] = 8'hAA;
ROM_MEM[1583] = 8'hBC;
ROM_MEM[1584] = 8'hD9;
ROM_MEM[1585] = 8'hAA;
ROM_MEM[1586] = 8'hA4;
ROM_MEM[1587] = 8'h50;
ROM_MEM[1588] = 8'hBA;
ROM_MEM[1589] = 8'hCC;
ROM_MEM[1590] = 8'h50;
ROM_MEM[1591] = 8'h8F;
ROM_MEM[1592] = 8'h1C;
ROM_MEM[1593] = 8'h62;
ROM_MEM[1594] = 8'hAF;
ROM_MEM[1595] = 8'h43;
ROM_MEM[1596] = 8'hDD;
ROM_MEM[1597] = 8'hCC;
ROM_MEM[1598] = 8'h89;
ROM_MEM[1599] = 8'h02;
ROM_MEM[1600] = 8'h7C;
ROM_MEM[1601] = 8'h66;
ROM_MEM[1602] = 8'h2E;
ROM_MEM[1603] = 8'h6E;
ROM_MEM[1604] = 8'h70;
ROM_MEM[1605] = 8'h25;
ROM_MEM[1606] = 8'h9E;
ROM_MEM[1607] = 8'h56;
ROM_MEM[1608] = 8'h69;
ROM_MEM[1609] = 8'hB8;
ROM_MEM[1610] = 8'hB6;
ROM_MEM[1611] = 8'hAC;
ROM_MEM[1612] = 8'h79;
ROM_MEM[1613] = 8'hE9;
ROM_MEM[1614] = 8'h98;
ROM_MEM[1615] = 8'hE1;
ROM_MEM[1616] = 8'hD9;
ROM_MEM[1617] = 8'h55;
ROM_MEM[1618] = 8'hEA;
ROM_MEM[1619] = 8'hE1;
ROM_MEM[1620] = 8'h73;
ROM_MEM[1621] = 8'h87;
ROM_MEM[1622] = 8'h67;
ROM_MEM[1623] = 8'h77;
ROM_MEM[1624] = 8'hB8;
ROM_MEM[1625] = 8'h59;
ROM_MEM[1626] = 8'h2E;
ROM_MEM[1627] = 8'h69;
ROM_MEM[1628] = 8'hAE;
ROM_MEM[1629] = 8'hD9;
ROM_MEM[1630] = 8'hE9;
ROM_MEM[1631] = 8'h61;
ROM_MEM[1632] = 8'h51;
ROM_MEM[1633] = 8'h67;
ROM_MEM[1634] = 8'hB8;
ROM_MEM[1635] = 8'hFE;
ROM_MEM[1636] = 8'hAA;
ROM_MEM[1637] = 8'h7A;
ROM_MEM[1638] = 8'h64;
ROM_MEM[1639] = 8'h93;
ROM_MEM[1640] = 8'hE5;
ROM_MEM[1641] = 8'hC4;
ROM_MEM[1642] = 8'hCE;
ROM_MEM[1643] = 8'h91;
ROM_MEM[1644] = 8'h9D;
ROM_MEM[1645] = 8'h89;
ROM_MEM[1646] = 8'h97;
ROM_MEM[1647] = 8'h93;
ROM_MEM[1648] = 8'hA2;
ROM_MEM[1649] = 8'hA4;
ROM_MEM[1650] = 8'h4E;
ROM_MEM[1651] = 8'h24;
ROM_MEM[1652] = 8'h5C;
ROM_MEM[1653] = 8'h76;
ROM_MEM[1654] = 8'h4E;
ROM_MEM[1655] = 8'h14;
ROM_MEM[1656] = 8'h59;
ROM_MEM[1657] = 8'h69;
ROM_MEM[1658] = 8'hE5;
ROM_MEM[1659] = 8'h38;
ROM_MEM[1660] = 8'hB5;
ROM_MEM[1661] = 8'h90;
ROM_MEM[1662] = 8'hD6;
ROM_MEM[1663] = 8'h94;
ROM_MEM[1664] = 8'h95;
ROM_MEM[1665] = 8'hE3;
ROM_MEM[1666] = 8'hD6;
ROM_MEM[1667] = 8'h4C;
ROM_MEM[1668] = 8'h16;
ROM_MEM[1669] = 8'hD3;
ROM_MEM[1670] = 8'h76;
ROM_MEM[1671] = 8'h8E;
ROM_MEM[1672] = 8'h5F;
ROM_MEM[1673] = 8'h23;
ROM_MEM[1674] = 8'h59;
ROM_MEM[1675] = 8'hCC;
ROM_MEM[1676] = 8'hD8;
ROM_MEM[1677] = 8'h39;
ROM_MEM[1678] = 8'h61;
ROM_MEM[1679] = 8'h2B;
ROM_MEM[1680] = 8'hCC;
ROM_MEM[1681] = 8'h51;
ROM_MEM[1682] = 8'h2B;
ROM_MEM[1683] = 8'hFB;
ROM_MEM[1684] = 8'hC4;
ROM_MEM[1685] = 8'h35;
ROM_MEM[1686] = 8'hB3;
ROM_MEM[1687] = 8'h66;
ROM_MEM[1688] = 8'hAD;
ROM_MEM[1689] = 8'hED;
ROM_MEM[1690] = 8'h95;
ROM_MEM[1691] = 8'hD6;
ROM_MEM[1692] = 8'h42;
ROM_MEM[1693] = 8'h56;
ROM_MEM[1694] = 8'h35;
ROM_MEM[1695] = 8'h8A;
ROM_MEM[1696] = 8'h57;
ROM_MEM[1697] = 8'h5E;
ROM_MEM[1698] = 8'h0A;
ROM_MEM[1699] = 8'h4B;
ROM_MEM[1700] = 8'hE5;
ROM_MEM[1701] = 8'hC8;
ROM_MEM[1702] = 8'h1E;
ROM_MEM[1703] = 8'h65;
ROM_MEM[1704] = 8'h36;
ROM_MEM[1705] = 8'h41;
ROM_MEM[1706] = 8'h13;
ROM_MEM[1707] = 8'h6D;
ROM_MEM[1708] = 8'hA5;
ROM_MEM[1709] = 8'h15;
ROM_MEM[1710] = 8'h89;
ROM_MEM[1711] = 8'hBB;
ROM_MEM[1712] = 8'h95;
ROM_MEM[1713] = 8'hB6;
ROM_MEM[1714] = 8'hEC;
ROM_MEM[1715] = 8'h92;
ROM_MEM[1716] = 8'h07;
ROM_MEM[1717] = 8'h91;
ROM_MEM[1718] = 8'hD6;
ROM_MEM[1719] = 8'h9A;
ROM_MEM[1720] = 8'h72;
ROM_MEM[1721] = 8'h42;
ROM_MEM[1722] = 8'h16;
ROM_MEM[1723] = 8'h54;
ROM_MEM[1724] = 8'h98;
ROM_MEM[1725] = 8'hB9;
ROM_MEM[1726] = 8'hD9;
ROM_MEM[1727] = 8'h7E;
ROM_MEM[1728] = 8'h80;
ROM_MEM[1729] = 8'h35;
ROM_MEM[1730] = 8'hA6;
ROM_MEM[1731] = 8'h8D;
ROM_MEM[1732] = 8'h8F;
ROM_MEM[1733] = 8'hA9;
ROM_MEM[1734] = 8'hCA;
ROM_MEM[1735] = 8'hC2;
ROM_MEM[1736] = 8'hEB;
ROM_MEM[1737] = 8'h2C;
ROM_MEM[1738] = 8'h21;
ROM_MEM[1739] = 8'hA6;
ROM_MEM[1740] = 8'hA9;
ROM_MEM[1741] = 8'hB4;
ROM_MEM[1742] = 8'h68;
ROM_MEM[1743] = 8'hB2;
ROM_MEM[1744] = 8'hE8;
ROM_MEM[1745] = 8'h14;
ROM_MEM[1746] = 8'hCE;
ROM_MEM[1747] = 8'hD3;
ROM_MEM[1748] = 8'h2D;
ROM_MEM[1749] = 8'hCE;
ROM_MEM[1750] = 8'hA2;
ROM_MEM[1751] = 8'h4A;
ROM_MEM[1752] = 8'h1E;
ROM_MEM[1753] = 8'h8B;
ROM_MEM[1754] = 8'h50;
ROM_MEM[1755] = 8'h5F;
ROM_MEM[1756] = 8'h83;
ROM_MEM[1757] = 8'hC9;
ROM_MEM[1758] = 8'h85;
ROM_MEM[1759] = 8'hA2;
ROM_MEM[1760] = 8'h2A;
ROM_MEM[1761] = 8'h96;
ROM_MEM[1762] = 8'h26;
ROM_MEM[1763] = 8'hA1;
ROM_MEM[1764] = 8'h14;
ROM_MEM[1765] = 8'h94;
ROM_MEM[1766] = 8'h0E;
ROM_MEM[1767] = 8'hB3;
ROM_MEM[1768] = 8'h1D;
ROM_MEM[1769] = 8'hEC;
ROM_MEM[1770] = 8'h9C;
ROM_MEM[1771] = 8'hCB;
ROM_MEM[1772] = 8'hDD;
ROM_MEM[1773] = 8'h2C;
ROM_MEM[1774] = 8'h96;
ROM_MEM[1775] = 8'h03;
ROM_MEM[1776] = 8'h12;
ROM_MEM[1777] = 8'h2F;
ROM_MEM[1778] = 8'h29;
ROM_MEM[1779] = 8'h40;
ROM_MEM[1780] = 8'h67;
ROM_MEM[1781] = 8'hCE;
ROM_MEM[1782] = 8'h8B;
ROM_MEM[1783] = 8'hCA;
ROM_MEM[1784] = 8'h42;
ROM_MEM[1785] = 8'hB9;
ROM_MEM[1786] = 8'hBB;
ROM_MEM[1787] = 8'h62;
ROM_MEM[1788] = 8'h2D;
ROM_MEM[1789] = 8'h32;
ROM_MEM[1790] = 8'h3B;
ROM_MEM[1791] = 8'h65;
ROM_MEM[1792] = 8'hF7;
ROM_MEM[1793] = 8'h98;
ROM_MEM[1794] = 8'hDD;
ROM_MEM[1795] = 8'hE8;
ROM_MEM[1796] = 8'hA0;
ROM_MEM[1797] = 8'h43;
ROM_MEM[1798] = 8'hC2;
ROM_MEM[1799] = 8'h72;
ROM_MEM[1800] = 8'h75;
ROM_MEM[1801] = 8'hE1;
ROM_MEM[1802] = 8'h92;
ROM_MEM[1803] = 8'h26;
ROM_MEM[1804] = 8'h5B;
ROM_MEM[1805] = 8'hF7;
ROM_MEM[1806] = 8'h58;
ROM_MEM[1807] = 8'h89;
ROM_MEM[1808] = 8'h1D;
ROM_MEM[1809] = 8'hD2;
ROM_MEM[1810] = 8'h58;
ROM_MEM[1811] = 8'hD5;
ROM_MEM[1812] = 8'h5C;
ROM_MEM[1813] = 8'h17;
ROM_MEM[1814] = 8'h60;
ROM_MEM[1815] = 8'h68;
ROM_MEM[1816] = 8'hA3;
ROM_MEM[1817] = 8'hC1;
ROM_MEM[1818] = 8'h14;
ROM_MEM[1819] = 8'h6A;
ROM_MEM[1820] = 8'h92;
ROM_MEM[1821] = 8'h11;
ROM_MEM[1822] = 8'h89;
ROM_MEM[1823] = 8'h07;
ROM_MEM[1824] = 8'h1D;
ROM_MEM[1825] = 8'h7C;
ROM_MEM[1826] = 8'h8A;
ROM_MEM[1827] = 8'h97;
ROM_MEM[1828] = 8'h24;
ROM_MEM[1829] = 8'h3A;
ROM_MEM[1830] = 8'h74;
ROM_MEM[1831] = 8'h74;
ROM_MEM[1832] = 8'hE5;
ROM_MEM[1833] = 8'hE1;
ROM_MEM[1834] = 8'hDE;
ROM_MEM[1835] = 8'h79;
ROM_MEM[1836] = 8'hD1;
ROM_MEM[1837] = 8'hB9;
ROM_MEM[1838] = 8'hA4;
ROM_MEM[1839] = 8'hBB;
ROM_MEM[1840] = 8'h7A;
ROM_MEM[1841] = 8'hEB;
ROM_MEM[1842] = 8'h43;
ROM_MEM[1843] = 8'h77;
ROM_MEM[1844] = 8'h97;
ROM_MEM[1845] = 8'h61;
ROM_MEM[1846] = 8'h66;
ROM_MEM[1847] = 8'hAD;
ROM_MEM[1848] = 8'h17;
ROM_MEM[1849] = 8'h3B;
ROM_MEM[1850] = 8'hB2;
ROM_MEM[1851] = 8'h17;
ROM_MEM[1852] = 8'h69;
ROM_MEM[1853] = 8'hCC;
ROM_MEM[1854] = 8'h69;
ROM_MEM[1855] = 8'h7C;
ROM_MEM[1856] = 8'h51;
ROM_MEM[1857] = 8'h1C;
ROM_MEM[1858] = 8'h21;
ROM_MEM[1859] = 8'h15;
ROM_MEM[1860] = 8'hF9;
ROM_MEM[1861] = 8'h08;
ROM_MEM[1862] = 8'h23;
ROM_MEM[1863] = 8'h8A;
ROM_MEM[1864] = 8'h69;
ROM_MEM[1865] = 8'h44;
ROM_MEM[1866] = 8'hED;
ROM_MEM[1867] = 8'h25;
ROM_MEM[1868] = 8'h0F;
ROM_MEM[1869] = 8'h2F;
ROM_MEM[1870] = 8'hEC;
ROM_MEM[1871] = 8'h1D;
ROM_MEM[1872] = 8'h8B;
ROM_MEM[1873] = 8'h82;
ROM_MEM[1874] = 8'h19;
ROM_MEM[1875] = 8'h85;
ROM_MEM[1876] = 8'h86;
ROM_MEM[1877] = 8'hBB;
ROM_MEM[1878] = 8'hDB;
ROM_MEM[1879] = 8'h0E;
ROM_MEM[1880] = 8'h41;
ROM_MEM[1881] = 8'hD3;
ROM_MEM[1882] = 8'hAA;
ROM_MEM[1883] = 8'h2E;
ROM_MEM[1884] = 8'h6A;
ROM_MEM[1885] = 8'h2B;
ROM_MEM[1886] = 8'h00;
ROM_MEM[1887] = 8'hA9;
ROM_MEM[1888] = 8'hB8;
ROM_MEM[1889] = 8'h34;
ROM_MEM[1890] = 8'hAE;
ROM_MEM[1891] = 8'h7A;
ROM_MEM[1892] = 8'h0F;
ROM_MEM[1893] = 8'h61;
ROM_MEM[1894] = 8'h8B;
ROM_MEM[1895] = 8'h73;
ROM_MEM[1896] = 8'hF8;
ROM_MEM[1897] = 8'h12;
ROM_MEM[1898] = 8'h9C;
ROM_MEM[1899] = 8'hA8;
ROM_MEM[1900] = 8'h2D;
ROM_MEM[1901] = 8'hF6;
ROM_MEM[1902] = 8'hE1;
ROM_MEM[1903] = 8'h87;
ROM_MEM[1904] = 8'h36;
ROM_MEM[1905] = 8'hE1;
ROM_MEM[1906] = 8'hF1;
ROM_MEM[1907] = 8'h38;
ROM_MEM[1908] = 8'h47;
ROM_MEM[1909] = 8'h18;
ROM_MEM[1910] = 8'hD9;
ROM_MEM[1911] = 8'h98;
ROM_MEM[1912] = 8'h2D;
ROM_MEM[1913] = 8'h66;
ROM_MEM[1914] = 8'h15;
ROM_MEM[1915] = 8'hB5;
ROM_MEM[1916] = 8'h69;
ROM_MEM[1917] = 8'h16;
ROM_MEM[1918] = 8'hCD;
ROM_MEM[1919] = 8'h88;
ROM_MEM[1920] = 8'h94;
ROM_MEM[1921] = 8'hB4;
ROM_MEM[1922] = 8'hE9;
ROM_MEM[1923] = 8'h5C;
ROM_MEM[1924] = 8'h58;
ROM_MEM[1925] = 8'hCC;
ROM_MEM[1926] = 8'hB1;
ROM_MEM[1927] = 8'h01;
ROM_MEM[1928] = 8'h1C;
ROM_MEM[1929] = 8'hB3;
ROM_MEM[1930] = 8'h38;
ROM_MEM[1931] = 8'h42;
ROM_MEM[1932] = 8'h53;
ROM_MEM[1933] = 8'hE2;
ROM_MEM[1934] = 8'hA1;
ROM_MEM[1935] = 8'h3E;
ROM_MEM[1936] = 8'hA9;
ROM_MEM[1937] = 8'hA8;
ROM_MEM[1938] = 8'h55;
ROM_MEM[1939] = 8'h6A;
ROM_MEM[1940] = 8'h98;
ROM_MEM[1941] = 8'hF1;
ROM_MEM[1942] = 8'hE4;
ROM_MEM[1943] = 8'hE0;
ROM_MEM[1944] = 8'h65;
ROM_MEM[1945] = 8'h4E;
ROM_MEM[1946] = 8'h9E;
ROM_MEM[1947] = 8'h6E;
ROM_MEM[1948] = 8'h8E;
ROM_MEM[1949] = 8'h04;
ROM_MEM[1950] = 8'h20;
ROM_MEM[1951] = 8'h84;
ROM_MEM[1952] = 8'h79;
ROM_MEM[1953] = 8'hE3;
ROM_MEM[1954] = 8'h9A;
ROM_MEM[1955] = 8'h16;
ROM_MEM[1956] = 8'h33;
ROM_MEM[1957] = 8'h97;
ROM_MEM[1958] = 8'hD2;
ROM_MEM[1959] = 8'h47;
ROM_MEM[1960] = 8'h4A;
ROM_MEM[1961] = 8'hA9;
ROM_MEM[1962] = 8'hC3;
ROM_MEM[1963] = 8'hCD;
ROM_MEM[1964] = 8'h82;
ROM_MEM[1965] = 8'h1C;
ROM_MEM[1966] = 8'hA9;
ROM_MEM[1967] = 8'hB8;
ROM_MEM[1968] = 8'hAE;
ROM_MEM[1969] = 8'hCA;
ROM_MEM[1970] = 8'h98;
ROM_MEM[1971] = 8'h74;
ROM_MEM[1972] = 8'hA4;
ROM_MEM[1973] = 8'h1C;
ROM_MEM[1974] = 8'hA6;
ROM_MEM[1975] = 8'h2B;
ROM_MEM[1976] = 8'h7D;
ROM_MEM[1977] = 8'hF2;
ROM_MEM[1978] = 8'h91;
ROM_MEM[1979] = 8'hB2;
ROM_MEM[1980] = 8'h9F;
ROM_MEM[1981] = 8'h9E;
ROM_MEM[1982] = 8'hB4;
ROM_MEM[1983] = 8'h9A;
ROM_MEM[1984] = 8'h43;
ROM_MEM[1985] = 8'hCE;
ROM_MEM[1986] = 8'h7E;
ROM_MEM[1987] = 8'h27;
ROM_MEM[1988] = 8'h4B;
ROM_MEM[1989] = 8'h1B;
ROM_MEM[1990] = 8'h0D;
ROM_MEM[1991] = 8'h25;
ROM_MEM[1992] = 8'hF9;
ROM_MEM[1993] = 8'hEB;
ROM_MEM[1994] = 8'h68;
ROM_MEM[1995] = 8'h69;
ROM_MEM[1996] = 8'h3A;
ROM_MEM[1997] = 8'h8C;
ROM_MEM[1998] = 8'h14;
ROM_MEM[1999] = 8'h76;
ROM_MEM[2000] = 8'h34;
ROM_MEM[2001] = 8'h6D;
ROM_MEM[2002] = 8'h6E;
ROM_MEM[2003] = 8'h73;
ROM_MEM[2004] = 8'h62;
ROM_MEM[2005] = 8'hB9;
ROM_MEM[2006] = 8'h91;
ROM_MEM[2007] = 8'hA0;
ROM_MEM[2008] = 8'h39;
ROM_MEM[2009] = 8'hCD;
ROM_MEM[2010] = 8'h8F;
ROM_MEM[2011] = 8'h71;
ROM_MEM[2012] = 8'h0B;
ROM_MEM[2013] = 8'hCB;
ROM_MEM[2014] = 8'hDB;
ROM_MEM[2015] = 8'hB4;
ROM_MEM[2016] = 8'h28;
ROM_MEM[2017] = 8'hBB;
ROM_MEM[2018] = 8'h1B;
ROM_MEM[2019] = 8'h4C;
ROM_MEM[2020] = 8'hAD;
ROM_MEM[2021] = 8'h3B;
ROM_MEM[2022] = 8'hD2;
ROM_MEM[2023] = 8'h62;
ROM_MEM[2024] = 8'h26;
ROM_MEM[2025] = 8'hA9;
ROM_MEM[2026] = 8'h2D;
ROM_MEM[2027] = 8'hDE;
ROM_MEM[2028] = 8'hCA;
ROM_MEM[2029] = 8'h8B;
ROM_MEM[2030] = 8'h9D;
ROM_MEM[2031] = 8'hA0;
ROM_MEM[2032] = 8'hD2;
ROM_MEM[2033] = 8'h26;
ROM_MEM[2034] = 8'hA3;
ROM_MEM[2035] = 8'hC8;
ROM_MEM[2036] = 8'hA9;
ROM_MEM[2037] = 8'hC5;
ROM_MEM[2038] = 8'h52;
ROM_MEM[2039] = 8'h1A;
ROM_MEM[2040] = 8'h97;
ROM_MEM[2041] = 8'hA2;
ROM_MEM[2042] = 8'h39;
ROM_MEM[2043] = 8'h17;
ROM_MEM[2044] = 8'h4D;
ROM_MEM[2045] = 8'h89;
ROM_MEM[2046] = 8'hF3;
ROM_MEM[2047] = 8'h00;
ROM_MEM[2048] = 8'h6E;
ROM_MEM[2049] = 8'h83;
ROM_MEM[2050] = 8'h29;
ROM_MEM[2051] = 8'h4E;
ROM_MEM[2052] = 8'h1F;
ROM_MEM[2053] = 8'h1C;
ROM_MEM[2054] = 8'h93;
ROM_MEM[2055] = 8'hBC;
ROM_MEM[2056] = 8'h23;
ROM_MEM[2057] = 8'h0D;
ROM_MEM[2058] = 8'h65;
ROM_MEM[2059] = 8'h5A;
ROM_MEM[2060] = 8'h4D;
ROM_MEM[2061] = 8'hF0;
ROM_MEM[2062] = 8'h8A;
ROM_MEM[2063] = 8'h72;
ROM_MEM[2064] = 8'hC4;
ROM_MEM[2065] = 8'h5A;
ROM_MEM[2066] = 8'h42;
ROM_MEM[2067] = 8'h70;
ROM_MEM[2068] = 8'hB5;
ROM_MEM[2069] = 8'hF5;
ROM_MEM[2070] = 8'hE2;
ROM_MEM[2071] = 8'h9A;
ROM_MEM[2072] = 8'hAB;
ROM_MEM[2073] = 8'hC4;
ROM_MEM[2074] = 8'hA3;
ROM_MEM[2075] = 8'hA6;
ROM_MEM[2076] = 8'h85;
ROM_MEM[2077] = 8'hCE;
ROM_MEM[2078] = 8'hBB;
ROM_MEM[2079] = 8'h9D;
ROM_MEM[2080] = 8'h87;
ROM_MEM[2081] = 8'hB3;
ROM_MEM[2082] = 8'h0E;
ROM_MEM[2083] = 8'hB2;
ROM_MEM[2084] = 8'hA4;
ROM_MEM[2085] = 8'h08;
ROM_MEM[2086] = 8'h2B;
ROM_MEM[2087] = 8'hDE;
ROM_MEM[2088] = 8'h76;
ROM_MEM[2089] = 8'h88;
ROM_MEM[2090] = 8'hAE;
ROM_MEM[2091] = 8'h7C;
ROM_MEM[2092] = 8'h74;
ROM_MEM[2093] = 8'h24;
ROM_MEM[2094] = 8'hF5;
ROM_MEM[2095] = 8'h22;
ROM_MEM[2096] = 8'h9A;
ROM_MEM[2097] = 8'h98;
ROM_MEM[2098] = 8'hA9;
ROM_MEM[2099] = 8'h16;
ROM_MEM[2100] = 8'h67;
ROM_MEM[2101] = 8'h0B;
ROM_MEM[2102] = 8'h6F;
ROM_MEM[2103] = 8'h72;
ROM_MEM[2104] = 8'hA6;
ROM_MEM[2105] = 8'h8A;
ROM_MEM[2106] = 8'hDD;
ROM_MEM[2107] = 8'h0D;
ROM_MEM[2108] = 8'hBC;
ROM_MEM[2109] = 8'h89;
ROM_MEM[2110] = 8'hD9;
ROM_MEM[2111] = 8'h0C;
ROM_MEM[2112] = 8'h71;
ROM_MEM[2113] = 8'h3F;
ROM_MEM[2114] = 8'h88;
ROM_MEM[2115] = 8'h26;
ROM_MEM[2116] = 8'h66;
ROM_MEM[2117] = 8'h2B;
ROM_MEM[2118] = 8'hC4;
ROM_MEM[2119] = 8'hF9;
ROM_MEM[2120] = 8'h20;
ROM_MEM[2121] = 8'h9A;
ROM_MEM[2122] = 8'hAC;
ROM_MEM[2123] = 8'h5D;
ROM_MEM[2124] = 8'hE3;
ROM_MEM[2125] = 8'hA4;
ROM_MEM[2126] = 8'h8B;
ROM_MEM[2127] = 8'h1C;
ROM_MEM[2128] = 8'hC6;
ROM_MEM[2129] = 8'hE2;
ROM_MEM[2130] = 8'h9C;
ROM_MEM[2131] = 8'hA7;
ROM_MEM[2132] = 8'h04;
ROM_MEM[2133] = 8'h20;
ROM_MEM[2134] = 8'hEA;
ROM_MEM[2135] = 8'h32;
ROM_MEM[2136] = 8'h01;
ROM_MEM[2137] = 8'h70;
ROM_MEM[2138] = 8'hDD;
ROM_MEM[2139] = 8'h0A;
ROM_MEM[2140] = 8'h09;
ROM_MEM[2141] = 8'h48;
ROM_MEM[2142] = 8'h52;
ROM_MEM[2143] = 8'h3D;
ROM_MEM[2144] = 8'h01;
ROM_MEM[2145] = 8'h45;
ROM_MEM[2146] = 8'hA7;
ROM_MEM[2147] = 8'h27;
ROM_MEM[2148] = 8'hB2;
ROM_MEM[2149] = 8'h8A;
ROM_MEM[2150] = 8'hCA;
ROM_MEM[2151] = 8'h40;
ROM_MEM[2152] = 8'h71;
ROM_MEM[2153] = 8'h5C;
ROM_MEM[2154] = 8'h88;
ROM_MEM[2155] = 8'h22;
ROM_MEM[2156] = 8'hAD;
ROM_MEM[2157] = 8'h4D;
ROM_MEM[2158] = 8'h24;
ROM_MEM[2159] = 8'hED;
ROM_MEM[2160] = 8'hC0;
ROM_MEM[2161] = 8'h73;
ROM_MEM[2162] = 8'hE8;
ROM_MEM[2163] = 8'h31;
ROM_MEM[2164] = 8'hA1;
ROM_MEM[2165] = 8'hB9;
ROM_MEM[2166] = 8'h0B;
ROM_MEM[2167] = 8'h6F;
ROM_MEM[2168] = 8'h2E;
ROM_MEM[2169] = 8'hBA;
ROM_MEM[2170] = 8'h8A;
ROM_MEM[2171] = 8'hC7;
ROM_MEM[2172] = 8'h1E;
ROM_MEM[2173] = 8'h7C;
ROM_MEM[2174] = 8'h86;
ROM_MEM[2175] = 8'h4C;
ROM_MEM[2176] = 8'h1D;
ROM_MEM[2177] = 8'h29;
ROM_MEM[2178] = 8'h7B;
ROM_MEM[2179] = 8'h88;
ROM_MEM[2180] = 8'h11;
ROM_MEM[2181] = 8'h67;
ROM_MEM[2182] = 8'hB8;
ROM_MEM[2183] = 8'h2C;
ROM_MEM[2184] = 8'hC9;
ROM_MEM[2185] = 8'h22;
ROM_MEM[2186] = 8'hEB;
ROM_MEM[2187] = 8'hBE;
ROM_MEM[2188] = 8'hD6;
ROM_MEM[2189] = 8'hD0;
ROM_MEM[2190] = 8'h3A;
ROM_MEM[2191] = 8'h8B;
ROM_MEM[2192] = 8'hAA;
ROM_MEM[2193] = 8'h6D;
ROM_MEM[2194] = 8'h5B;
ROM_MEM[2195] = 8'h8A;
ROM_MEM[2196] = 8'hEB;
ROM_MEM[2197] = 8'h2C;
ROM_MEM[2198] = 8'hBA;
ROM_MEM[2199] = 8'hD6;
ROM_MEM[2200] = 8'h29;
ROM_MEM[2201] = 8'h29;
ROM_MEM[2202] = 8'h4A;
ROM_MEM[2203] = 8'hD2;
ROM_MEM[2204] = 8'hC4;
ROM_MEM[2205] = 8'h36;
ROM_MEM[2206] = 8'hC2;
ROM_MEM[2207] = 8'h34;
ROM_MEM[2208] = 8'hB9;
ROM_MEM[2209] = 8'hA5;
ROM_MEM[2210] = 8'h33;
ROM_MEM[2211] = 8'h6A;
ROM_MEM[2212] = 8'h51;
ROM_MEM[2213] = 8'h92;
ROM_MEM[2214] = 8'h90;
ROM_MEM[2215] = 8'hD4;
ROM_MEM[2216] = 8'hD0;
ROM_MEM[2217] = 8'h80;
ROM_MEM[2218] = 8'h4E;
ROM_MEM[2219] = 8'h89;
ROM_MEM[2220] = 8'h12;
ROM_MEM[2221] = 8'hD0;
ROM_MEM[2222] = 8'hA5;
ROM_MEM[2223] = 8'h78;
ROM_MEM[2224] = 8'h13;
ROM_MEM[2225] = 8'hA6;
ROM_MEM[2226] = 8'h16;
ROM_MEM[2227] = 8'hB6;
ROM_MEM[2228] = 8'h88;
ROM_MEM[2229] = 8'hD8;
ROM_MEM[2230] = 8'h87;
ROM_MEM[2231] = 8'h1E;
ROM_MEM[2232] = 8'h7D;
ROM_MEM[2233] = 8'h12;
ROM_MEM[2234] = 8'h3C;
ROM_MEM[2235] = 8'hAD;
ROM_MEM[2236] = 8'h1C;
ROM_MEM[2237] = 8'h7A;
ROM_MEM[2238] = 8'hE4;
ROM_MEM[2239] = 8'h34;
ROM_MEM[2240] = 8'h9E;
ROM_MEM[2241] = 8'h88;
ROM_MEM[2242] = 8'h77;
ROM_MEM[2243] = 8'hA8;
ROM_MEM[2244] = 8'hE1;
ROM_MEM[2245] = 8'hCD;
ROM_MEM[2246] = 8'hAD;
ROM_MEM[2247] = 8'hB4;
ROM_MEM[2248] = 8'hED;
ROM_MEM[2249] = 8'hA1;
ROM_MEM[2250] = 8'h46;
ROM_MEM[2251] = 8'hF3;
ROM_MEM[2252] = 8'h4C;
ROM_MEM[2253] = 8'hB5;
ROM_MEM[2254] = 8'hB2;
ROM_MEM[2255] = 8'h84;
ROM_MEM[2256] = 8'hEE;
ROM_MEM[2257] = 8'hC5;
ROM_MEM[2258] = 8'h9C;
ROM_MEM[2259] = 8'hAC;
ROM_MEM[2260] = 8'hA2;
ROM_MEM[2261] = 8'h12;
ROM_MEM[2262] = 8'hBA;
ROM_MEM[2263] = 8'h69;
ROM_MEM[2264] = 8'h8A;
ROM_MEM[2265] = 8'hF2;
ROM_MEM[2266] = 8'h36;
ROM_MEM[2267] = 8'hF3;
ROM_MEM[2268] = 8'h00;
ROM_MEM[2269] = 8'h8B;
ROM_MEM[2270] = 8'hAE;
ROM_MEM[2271] = 8'hE2;
ROM_MEM[2272] = 8'h69;
ROM_MEM[2273] = 8'h88;
ROM_MEM[2274] = 8'h32;
ROM_MEM[2275] = 8'hCC;
ROM_MEM[2276] = 8'h3C;
ROM_MEM[2277] = 8'h27;
ROM_MEM[2278] = 8'h9F;
ROM_MEM[2279] = 8'hA4;
ROM_MEM[2280] = 8'h26;
ROM_MEM[2281] = 8'h0D;
ROM_MEM[2282] = 8'hF1;
ROM_MEM[2283] = 8'h34;
ROM_MEM[2284] = 8'h7D;
ROM_MEM[2285] = 8'hC2;
ROM_MEM[2286] = 8'h56;
ROM_MEM[2287] = 8'h38;
ROM_MEM[2288] = 8'hB1;
ROM_MEM[2289] = 8'hC3;
ROM_MEM[2290] = 8'hF2;
ROM_MEM[2291] = 8'hF1;
ROM_MEM[2292] = 8'h6B;
ROM_MEM[2293] = 8'hA6;
ROM_MEM[2294] = 8'hE0;
ROM_MEM[2295] = 8'h2E;
ROM_MEM[2296] = 8'h2B;
ROM_MEM[2297] = 8'h25;
ROM_MEM[2298] = 8'h19;
ROM_MEM[2299] = 8'hCA;
ROM_MEM[2300] = 8'h51;
ROM_MEM[2301] = 8'hC3;
ROM_MEM[2302] = 8'h2C;
ROM_MEM[2303] = 8'h13;
ROM_MEM[2304] = 8'hC0;
ROM_MEM[2305] = 8'h1A;
ROM_MEM[2306] = 8'h37;
ROM_MEM[2307] = 8'h04;
ROM_MEM[2308] = 8'h38;
ROM_MEM[2309] = 8'hE9;
ROM_MEM[2310] = 8'h21;
ROM_MEM[2311] = 8'h80;
ROM_MEM[2312] = 8'hA2;
ROM_MEM[2313] = 8'h5D;
ROM_MEM[2314] = 8'h11;
ROM_MEM[2315] = 8'h10;
ROM_MEM[2316] = 8'h99;
ROM_MEM[2317] = 8'h39;
ROM_MEM[2318] = 8'h02;
ROM_MEM[2319] = 8'hA8;
ROM_MEM[2320] = 8'hC8;
ROM_MEM[2321] = 8'h54;
ROM_MEM[2322] = 8'h69;
ROM_MEM[2323] = 8'h26;
ROM_MEM[2324] = 8'h62;
ROM_MEM[2325] = 8'h9E;
ROM_MEM[2326] = 8'h55;
ROM_MEM[2327] = 8'h67;
ROM_MEM[2328] = 8'h24;
ROM_MEM[2329] = 8'h75;
ROM_MEM[2330] = 8'hBB;
ROM_MEM[2331] = 8'hAB;
ROM_MEM[2332] = 8'h99;
ROM_MEM[2333] = 8'hAD;
ROM_MEM[2334] = 8'h11;
ROM_MEM[2335] = 8'h17;
ROM_MEM[2336] = 8'h27;
ROM_MEM[2337] = 8'h89;
ROM_MEM[2338] = 8'h91;
ROM_MEM[2339] = 8'h51;
ROM_MEM[2340] = 8'h56;
ROM_MEM[2341] = 8'h92;
ROM_MEM[2342] = 8'hA3;
ROM_MEM[2343] = 8'h37;
ROM_MEM[2344] = 8'h59;
ROM_MEM[2345] = 8'hC4;
ROM_MEM[2346] = 8'h3E;
ROM_MEM[2347] = 8'h61;
ROM_MEM[2348] = 8'hF6;
ROM_MEM[2349] = 8'hB1;
ROM_MEM[2350] = 8'hA4;
ROM_MEM[2351] = 8'h5E;
ROM_MEM[2352] = 8'hF7;
ROM_MEM[2353] = 8'hF8;
ROM_MEM[2354] = 8'hD5;
ROM_MEM[2355] = 8'hFA;
ROM_MEM[2356] = 8'h38;
ROM_MEM[2357] = 8'hF3;
ROM_MEM[2358] = 8'hDC;
ROM_MEM[2359] = 8'hE3;
ROM_MEM[2360] = 8'h25;
ROM_MEM[2361] = 8'h97;
ROM_MEM[2362] = 8'hC3;
ROM_MEM[2363] = 8'h1C;
ROM_MEM[2364] = 8'h53;
ROM_MEM[2365] = 8'h8F;
ROM_MEM[2366] = 8'h97;
ROM_MEM[2367] = 8'h7D;
ROM_MEM[2368] = 8'h0E;
ROM_MEM[2369] = 8'h93;
ROM_MEM[2370] = 8'h4F;
ROM_MEM[2371] = 8'h3D;
ROM_MEM[2372] = 8'h5E;
ROM_MEM[2373] = 8'h76;
ROM_MEM[2374] = 8'h39;
ROM_MEM[2375] = 8'h42;
ROM_MEM[2376] = 8'h3A;
ROM_MEM[2377] = 8'hED;
ROM_MEM[2378] = 8'h78;
ROM_MEM[2379] = 8'hC9;
ROM_MEM[2380] = 8'h55;
ROM_MEM[2381] = 8'h33;
ROM_MEM[2382] = 8'hFB;
ROM_MEM[2383] = 8'hDC;
ROM_MEM[2384] = 8'hE5;
ROM_MEM[2385] = 8'hC7;
ROM_MEM[2386] = 8'h50;
ROM_MEM[2387] = 8'h4D;
ROM_MEM[2388] = 8'h1C;
ROM_MEM[2389] = 8'h57;
ROM_MEM[2390] = 8'h47;
ROM_MEM[2391] = 8'h10;
ROM_MEM[2392] = 8'h5A;
ROM_MEM[2393] = 8'h27;
ROM_MEM[2394] = 8'h4A;
ROM_MEM[2395] = 8'h4C;
ROM_MEM[2396] = 8'h6B;
ROM_MEM[2397] = 8'h61;
ROM_MEM[2398] = 8'h38;
ROM_MEM[2399] = 8'hE9;
ROM_MEM[2400] = 8'hE0;
ROM_MEM[2401] = 8'h55;
ROM_MEM[2402] = 8'hB7;
ROM_MEM[2403] = 8'hC4;
ROM_MEM[2404] = 8'h61;
ROM_MEM[2405] = 8'h74;
ROM_MEM[2406] = 8'h82;
ROM_MEM[2407] = 8'h64;
ROM_MEM[2408] = 8'h99;
ROM_MEM[2409] = 8'h94;
ROM_MEM[2410] = 8'h87;
ROM_MEM[2411] = 8'h9B;
ROM_MEM[2412] = 8'h06;
ROM_MEM[2413] = 8'h56;
ROM_MEM[2414] = 8'h71;
ROM_MEM[2415] = 8'h42;
ROM_MEM[2416] = 8'hE5;
ROM_MEM[2417] = 8'hCB;
ROM_MEM[2418] = 8'h04;
ROM_MEM[2419] = 8'hA9;
ROM_MEM[2420] = 8'h25;
ROM_MEM[2421] = 8'h0D;
ROM_MEM[2422] = 8'h8D;
ROM_MEM[2423] = 8'h2F;
ROM_MEM[2424] = 8'hED;
ROM_MEM[2425] = 8'hA8;
ROM_MEM[2426] = 8'h9E;
ROM_MEM[2427] = 8'h26;
ROM_MEM[2428] = 8'hF4;
ROM_MEM[2429] = 8'h21;
ROM_MEM[2430] = 8'h76;
ROM_MEM[2431] = 8'h09;
ROM_MEM[2432] = 8'h85;
ROM_MEM[2433] = 8'h5D;
ROM_MEM[2434] = 8'h06;
ROM_MEM[2435] = 8'hA8;
ROM_MEM[2436] = 8'h9C;
ROM_MEM[2437] = 8'hCA;
ROM_MEM[2438] = 8'h00;
ROM_MEM[2439] = 8'hE1;
ROM_MEM[2440] = 8'hCB;
ROM_MEM[2441] = 8'h19;
ROM_MEM[2442] = 8'hA0;
ROM_MEM[2443] = 8'h7C;
ROM_MEM[2444] = 8'h28;
ROM_MEM[2445] = 8'h03;
ROM_MEM[2446] = 8'h44;
ROM_MEM[2447] = 8'h30;
ROM_MEM[2448] = 8'h27;
ROM_MEM[2449] = 8'h00;
ROM_MEM[2450] = 8'hCB;
ROM_MEM[2451] = 8'h69;
ROM_MEM[2452] = 8'h6E;
ROM_MEM[2453] = 8'hCE;
ROM_MEM[2454] = 8'h3A;
ROM_MEM[2455] = 8'h94;
ROM_MEM[2456] = 8'h2D;
ROM_MEM[2457] = 8'h9D;
ROM_MEM[2458] = 8'hA6;
ROM_MEM[2459] = 8'h39;
ROM_MEM[2460] = 8'h86;
ROM_MEM[2461] = 8'h30;
ROM_MEM[2462] = 8'hB5;
ROM_MEM[2463] = 8'h48;
ROM_MEM[2464] = 8'h9D;
ROM_MEM[2465] = 8'hA6;
ROM_MEM[2466] = 8'h10;
ROM_MEM[2467] = 8'h3C;
ROM_MEM[2468] = 8'h48;
ROM_MEM[2469] = 8'hBB;
ROM_MEM[2470] = 8'h4E;
ROM_MEM[2471] = 8'h9A;
ROM_MEM[2472] = 8'h9C;
ROM_MEM[2473] = 8'hCF;
ROM_MEM[2474] = 8'h14;
ROM_MEM[2475] = 8'hAD;
ROM_MEM[2476] = 8'h26;
ROM_MEM[2477] = 8'h61;
ROM_MEM[2478] = 8'h0E;
ROM_MEM[2479] = 8'hB9;
ROM_MEM[2480] = 8'h95;
ROM_MEM[2481] = 8'h24;
ROM_MEM[2482] = 8'h9B;
ROM_MEM[2483] = 8'hB8;
ROM_MEM[2484] = 8'h25;
ROM_MEM[2485] = 8'h98;
ROM_MEM[2486] = 8'h76;
ROM_MEM[2487] = 8'h61;
ROM_MEM[2488] = 8'h4B;
ROM_MEM[2489] = 8'hEA;
ROM_MEM[2490] = 8'hD6;
ROM_MEM[2491] = 8'h28;
ROM_MEM[2492] = 8'h2B;
ROM_MEM[2493] = 8'h54;
ROM_MEM[2494] = 8'hD4;
ROM_MEM[2495] = 8'h29;
ROM_MEM[2496] = 8'h01;
ROM_MEM[2497] = 8'hB4;
ROM_MEM[2498] = 8'h2B;
ROM_MEM[2499] = 8'h47;
ROM_MEM[2500] = 8'h80;
ROM_MEM[2501] = 8'h93;
ROM_MEM[2502] = 8'hE9;
ROM_MEM[2503] = 8'h08;
ROM_MEM[2504] = 8'hF0;
ROM_MEM[2505] = 8'h22;
ROM_MEM[2506] = 8'h1D;
ROM_MEM[2507] = 8'h18;
ROM_MEM[2508] = 8'h50;
ROM_MEM[2509] = 8'h82;
ROM_MEM[2510] = 8'h33;
ROM_MEM[2511] = 8'h01;
ROM_MEM[2512] = 8'h62;
ROM_MEM[2513] = 8'h0E;
ROM_MEM[2514] = 8'h79;
ROM_MEM[2515] = 8'h93;
ROM_MEM[2516] = 8'hE9;
ROM_MEM[2517] = 8'h08;
ROM_MEM[2518] = 8'h04;
ROM_MEM[2519] = 8'h68;
ROM_MEM[2520] = 8'hCC;
ROM_MEM[2521] = 8'h9A;
ROM_MEM[2522] = 8'h01;
ROM_MEM[2523] = 8'h9D;
ROM_MEM[2524] = 8'h68;
ROM_MEM[2525] = 8'h33;
ROM_MEM[2526] = 8'hA0;
ROM_MEM[2527] = 8'h61;
ROM_MEM[2528] = 8'h6B;
ROM_MEM[2529] = 8'h05;
ROM_MEM[2530] = 8'h74;
ROM_MEM[2531] = 8'hA4;
ROM_MEM[2532] = 8'h2D;
ROM_MEM[2533] = 8'h80;
ROM_MEM[2534] = 8'hC4;
ROM_MEM[2535] = 8'hEB;
ROM_MEM[2536] = 8'h14;
ROM_MEM[2537] = 8'h50;
ROM_MEM[2538] = 8'h68;
ROM_MEM[2539] = 8'h8C;
ROM_MEM[2540] = 8'h02;
ROM_MEM[2541] = 8'h1A;
ROM_MEM[2542] = 8'h95;
ROM_MEM[2543] = 8'h56;
ROM_MEM[2544] = 8'h40;
ROM_MEM[2545] = 8'hE3;
ROM_MEM[2546] = 8'hD2;
ROM_MEM[2547] = 8'h0A;
ROM_MEM[2548] = 8'h28;
ROM_MEM[2549] = 8'hA4;
ROM_MEM[2550] = 8'h46;
ROM_MEM[2551] = 8'h01;
ROM_MEM[2552] = 8'h95;
ROM_MEM[2553] = 8'hD8;
ROM_MEM[2554] = 8'h18;
ROM_MEM[2555] = 8'hA0;
ROM_MEM[2556] = 8'h52;
ROM_MEM[2557] = 8'h5B;
ROM_MEM[2558] = 8'h07;
ROM_MEM[2559] = 8'h34;
ROM_MEM[2560] = 8'h2A;
ROM_MEM[2561] = 8'h63;
ROM_MEM[2562] = 8'h80;
ROM_MEM[2563] = 8'h46;
ROM_MEM[2564] = 8'hB4;
ROM_MEM[2565] = 8'h0D;
ROM_MEM[2566] = 8'h90;
ROM_MEM[2567] = 8'h59;
ROM_MEM[2568] = 8'hAC;
ROM_MEM[2569] = 8'h01;
ROM_MEM[2570] = 8'h1A;
ROM_MEM[2571] = 8'h91;
ROM_MEM[2572] = 8'h32;
ROM_MEM[2573] = 8'h40;
ROM_MEM[2574] = 8'h67;
ROM_MEM[2575] = 8'hDC;
ROM_MEM[2576] = 8'h06;
ROM_MEM[2577] = 8'h68;
ROM_MEM[2578] = 8'hC8;
ROM_MEM[2579] = 8'h5A;
ROM_MEM[2580] = 8'h01;
ROM_MEM[2581] = 8'h15;
ROM_MEM[2582] = 8'hE5;
ROM_MEM[2583] = 8'h18;
ROM_MEM[2584] = 8'hA0;
ROM_MEM[2585] = 8'h51;
ROM_MEM[2586] = 8'h69;
ROM_MEM[2587] = 8'h05;
ROM_MEM[2588] = 8'h14;
ROM_MEM[2589] = 8'h56;
ROM_MEM[2590] = 8'h6B;
ROM_MEM[2591] = 8'h80;
ROM_MEM[2592] = 8'h42;
ROM_MEM[2593] = 8'h6B;
ROM_MEM[2594] = 8'h14;
ROM_MEM[2595] = 8'h50;
ROM_MEM[2596] = 8'h48;
ROM_MEM[2597] = 8'h8E;
ROM_MEM[2598] = 8'h01;
ROM_MEM[2599] = 8'h1A;
ROM_MEM[2600] = 8'hB5;
ROM_MEM[2601] = 8'h51;
ROM_MEM[2602] = 8'h40;
ROM_MEM[2603] = 8'hA5;
ROM_MEM[2604] = 8'h36;
ROM_MEM[2605] = 8'h0A;
ROM_MEM[2606] = 8'hA8;
ROM_MEM[2607] = 8'hD4;
ROM_MEM[2608] = 8'h56;
ROM_MEM[2609] = 8'h01;
ROM_MEM[2610] = 8'h99;
ROM_MEM[2611] = 8'hE7;
ROM_MEM[2612] = 8'h2A;
ROM_MEM[2613] = 8'hA0;
ROM_MEM[2614] = 8'hD0;
ROM_MEM[2615] = 8'h18;
ROM_MEM[2616] = 8'h01;
ROM_MEM[2617] = 8'h74;
ROM_MEM[2618] = 8'h6C;
ROM_MEM[2619] = 8'h2D;
ROM_MEM[2620] = 8'h80;
ROM_MEM[2621] = 8'hCE;
ROM_MEM[2622] = 8'hA4;
ROM_MEM[2623] = 8'h04;
ROM_MEM[2624] = 8'h50;
ROM_MEM[2625] = 8'h69;
ROM_MEM[2626] = 8'h34;
ROM_MEM[2627] = 8'h03;
ROM_MEM[2628] = 8'h1A;
ROM_MEM[2629] = 8'hF1;
ROM_MEM[2630] = 8'h66;
ROM_MEM[2631] = 8'h40;
ROM_MEM[2632] = 8'hA1;
ROM_MEM[2633] = 8'h35;
ROM_MEM[2634] = 8'h0C;
ROM_MEM[2635] = 8'hA8;
ROM_MEM[2636] = 8'h34;
ROM_MEM[2637] = 8'h86;
ROM_MEM[2638] = 8'h01;
ROM_MEM[2639] = 8'h8D;
ROM_MEM[2640] = 8'h69;
ROM_MEM[2641] = 8'h31;
ROM_MEM[2642] = 8'hA0;
ROM_MEM[2643] = 8'h31;
ROM_MEM[2644] = 8'hC9;
ROM_MEM[2645] = 8'h07;
ROM_MEM[2646] = 8'h54;
ROM_MEM[2647] = 8'h94;
ROM_MEM[2648] = 8'h63;
ROM_MEM[2649] = 8'hC6;
ROM_MEM[2650] = 8'hE9;
ROM_MEM[2651] = 8'h84;
ROM_MEM[2652] = 8'h35;
ROM_MEM[2653] = 8'hBA;
ROM_MEM[2654] = 8'hCC;
ROM_MEM[2655] = 8'h06;
ROM_MEM[2656] = 8'hB9;
ROM_MEM[2657] = 8'h73;
ROM_MEM[2658] = 8'h21;
ROM_MEM[2659] = 8'h1F;
ROM_MEM[2660] = 8'h8F;
ROM_MEM[2661] = 8'h33;
ROM_MEM[2662] = 8'hD8;
ROM_MEM[2663] = 8'hE1;
ROM_MEM[2664] = 8'h8C;
ROM_MEM[2665] = 8'h6C;
ROM_MEM[2666] = 8'h33;
ROM_MEM[2667] = 8'hCA;
ROM_MEM[2668] = 8'hA1;
ROM_MEM[2669] = 8'hAA;
ROM_MEM[2670] = 8'hD1;
ROM_MEM[2671] = 8'hC8;
ROM_MEM[2672] = 8'hCB;
ROM_MEM[2673] = 8'hA6;
ROM_MEM[2674] = 8'h87;
ROM_MEM[2675] = 8'h6A;
ROM_MEM[2676] = 8'h23;
ROM_MEM[2677] = 8'hCD;
ROM_MEM[2678] = 8'hC7;
ROM_MEM[2679] = 8'hED;
ROM_MEM[2680] = 8'h1C;
ROM_MEM[2681] = 8'hB2;
ROM_MEM[2682] = 8'hB6;
ROM_MEM[2683] = 8'hB4;
ROM_MEM[2684] = 8'hAC;
ROM_MEM[2685] = 8'h72;
ROM_MEM[2686] = 8'h7C;
ROM_MEM[2687] = 8'h88;
ROM_MEM[2688] = 8'h1A;
ROM_MEM[2689] = 8'hD6;
ROM_MEM[2690] = 8'hBA;
ROM_MEM[2691] = 8'hCA;
ROM_MEM[2692] = 8'hEE;
ROM_MEM[2693] = 8'hC1;
ROM_MEM[2694] = 8'h4B;
ROM_MEM[2695] = 8'h3E;
ROM_MEM[2696] = 8'hAD;
ROM_MEM[2697] = 8'h68;
ROM_MEM[2698] = 8'hC7;
ROM_MEM[2699] = 8'h07;
ROM_MEM[2700] = 8'h2B;
ROM_MEM[2701] = 8'hF9;
ROM_MEM[2702] = 8'h25;
ROM_MEM[2703] = 8'hBB;
ROM_MEM[2704] = 8'hA4;
ROM_MEM[2705] = 8'h1C;
ROM_MEM[2706] = 8'hAC;
ROM_MEM[2707] = 8'hE4;
ROM_MEM[2708] = 8'hD5;
ROM_MEM[2709] = 8'hCC;
ROM_MEM[2710] = 8'h94;
ROM_MEM[2711] = 8'h7B;
ROM_MEM[2712] = 8'hB0;
ROM_MEM[2713] = 8'h5C;
ROM_MEM[2714] = 8'h47;
ROM_MEM[2715] = 8'hBA;
ROM_MEM[2716] = 8'h42;
ROM_MEM[2717] = 8'hE9;
ROM_MEM[2718] = 8'hC1;
ROM_MEM[2719] = 8'h72;
ROM_MEM[2720] = 8'h1B;
ROM_MEM[2721] = 8'hAD;
ROM_MEM[2722] = 8'h0A;
ROM_MEM[2723] = 8'h25;
ROM_MEM[2724] = 8'h07;
ROM_MEM[2725] = 8'h2B;
ROM_MEM[2726] = 8'h73;
ROM_MEM[2727] = 8'h2C;
ROM_MEM[2728] = 8'hBA;
ROM_MEM[2729] = 8'h15;
ROM_MEM[2730] = 8'h0F;
ROM_MEM[2731] = 8'h2C;
ROM_MEM[2732] = 8'hE7;
ROM_MEM[2733] = 8'h51;
ROM_MEM[2734] = 8'hAB;
ROM_MEM[2735] = 8'h50;
ROM_MEM[2736] = 8'hB4;
ROM_MEM[2737] = 8'hA8;
ROM_MEM[2738] = 8'h54;
ROM_MEM[2739] = 8'h43;
ROM_MEM[2740] = 8'h63;
ROM_MEM[2741] = 8'h59;
ROM_MEM[2742] = 8'hF5;
ROM_MEM[2743] = 8'hA1;
ROM_MEM[2744] = 8'h52;
ROM_MEM[2745] = 8'h71;
ROM_MEM[2746] = 8'hF5;
ROM_MEM[2747] = 8'h53;
ROM_MEM[2748] = 8'h27;
ROM_MEM[2749] = 8'h87;
ROM_MEM[2750] = 8'h4E;
ROM_MEM[2751] = 8'h29;
ROM_MEM[2752] = 8'hD5;
ROM_MEM[2753] = 8'hC6;
ROM_MEM[2754] = 8'hEC;
ROM_MEM[2755] = 8'h1C;
ROM_MEM[2756] = 8'h3C;
ROM_MEM[2757] = 8'h87;
ROM_MEM[2758] = 8'h11;
ROM_MEM[2759] = 8'hCD;
ROM_MEM[2760] = 8'hB4;
ROM_MEM[2761] = 8'h7D;
ROM_MEM[2762] = 8'hD0;
ROM_MEM[2763] = 8'hEC;
ROM_MEM[2764] = 8'hC6;
ROM_MEM[2765] = 8'hD1;
ROM_MEM[2766] = 8'hC3;
ROM_MEM[2767] = 8'hCE;
ROM_MEM[2768] = 8'h41;
ROM_MEM[2769] = 8'h8B;
ROM_MEM[2770] = 8'h7D;
ROM_MEM[2771] = 8'h26;
ROM_MEM[2772] = 8'hCB;
ROM_MEM[2773] = 8'hA4;
ROM_MEM[2774] = 8'h07;
ROM_MEM[2775] = 8'hCD;
ROM_MEM[2776] = 8'h7E;
ROM_MEM[2777] = 8'h85;
ROM_MEM[2778] = 8'h2C;
ROM_MEM[2779] = 8'h16;
ROM_MEM[2780] = 8'h1F;
ROM_MEM[2781] = 8'h24;
ROM_MEM[2782] = 8'hFB;
ROM_MEM[2783] = 8'h56;
ROM_MEM[2784] = 8'h96;
ROM_MEM[2785] = 8'h9A;
ROM_MEM[2786] = 8'h7D;
ROM_MEM[2787] = 8'hD0;
ROM_MEM[2788] = 8'h64;
ROM_MEM[2789] = 8'h5B;
ROM_MEM[2790] = 8'h44;
ROM_MEM[2791] = 8'hAB;
ROM_MEM[2792] = 8'hF1;
ROM_MEM[2793] = 8'h42;
ROM_MEM[2794] = 8'h93;
ROM_MEM[2795] = 8'h6B;
ROM_MEM[2796] = 8'h61;
ROM_MEM[2797] = 8'hED;
ROM_MEM[2798] = 8'h25;
ROM_MEM[2799] = 8'h03;
ROM_MEM[2800] = 8'h8D;
ROM_MEM[2801] = 8'hA1;
ROM_MEM[2802] = 8'h84;
ROM_MEM[2803] = 8'hBC;
ROM_MEM[2804] = 8'h1B;
ROM_MEM[2805] = 8'h2F;
ROM_MEM[2806] = 8'h2C;
ROM_MEM[2807] = 8'hB9;
ROM_MEM[2808] = 8'h36;
ROM_MEM[2809] = 8'h96;
ROM_MEM[2810] = 8'h68;
ROM_MEM[2811] = 8'h32;
ROM_MEM[2812] = 8'hF0;
ROM_MEM[2813] = 8'hAC;
ROM_MEM[2814] = 8'h4F;
ROM_MEM[2815] = 8'hC8;
ROM_MEM[2816] = 8'h62;
ROM_MEM[2817] = 8'h49;
ROM_MEM[2818] = 8'h23;
ROM_MEM[2819] = 8'h92;
ROM_MEM[2820] = 8'h1B;
ROM_MEM[2821] = 8'h03;
ROM_MEM[2822] = 8'h8B;
ROM_MEM[2823] = 8'hBA;
ROM_MEM[2824] = 8'h85;
ROM_MEM[2825] = 8'h8A;
ROM_MEM[2826] = 8'h6E;
ROM_MEM[2827] = 8'h15;
ROM_MEM[2828] = 8'hCD;
ROM_MEM[2829] = 8'h9A;
ROM_MEM[2830] = 8'h25;
ROM_MEM[2831] = 8'h26;
ROM_MEM[2832] = 8'hB2;
ROM_MEM[2833] = 8'h09;
ROM_MEM[2834] = 8'h0A;
ROM_MEM[2835] = 8'hB7;
ROM_MEM[2836] = 8'h1B;
ROM_MEM[2837] = 8'hB8;
ROM_MEM[2838] = 8'h48;
ROM_MEM[2839] = 8'hBB;
ROM_MEM[2840] = 8'h39;
ROM_MEM[2841] = 8'hCC;
ROM_MEM[2842] = 8'h8E;
ROM_MEM[2843] = 8'h93;
ROM_MEM[2844] = 8'h83;
ROM_MEM[2845] = 8'hDC;
ROM_MEM[2846] = 8'hA0;
ROM_MEM[2847] = 8'hF0;
ROM_MEM[2848] = 8'h24;
ROM_MEM[2849] = 8'hC6;
ROM_MEM[2850] = 8'hF0;
ROM_MEM[2851] = 8'h7E;
ROM_MEM[2852] = 8'h8D;
ROM_MEM[2853] = 8'hCC;
ROM_MEM[2854] = 8'h9B;
ROM_MEM[2855] = 8'h18;
ROM_MEM[2856] = 8'hCF;
ROM_MEM[2857] = 8'hCB;
ROM_MEM[2858] = 8'h49;
ROM_MEM[2859] = 8'h36;
ROM_MEM[2860] = 8'h4F;
ROM_MEM[2861] = 8'h66;
ROM_MEM[2862] = 8'hE2;
ROM_MEM[2863] = 8'hC0;
ROM_MEM[2864] = 8'hA7;
ROM_MEM[2865] = 8'h4C;
ROM_MEM[2866] = 8'hDC;
ROM_MEM[2867] = 8'hE9;
ROM_MEM[2868] = 8'h03;
ROM_MEM[2869] = 8'h4A;
ROM_MEM[2870] = 8'h7E;
ROM_MEM[2871] = 8'hC9;
ROM_MEM[2872] = 8'h6D;
ROM_MEM[2873] = 8'hAD;
ROM_MEM[2874] = 8'h46;
ROM_MEM[2875] = 8'hA7;
ROM_MEM[2876] = 8'h5C;
ROM_MEM[2877] = 8'hED;
ROM_MEM[2878] = 8'h8C;
ROM_MEM[2879] = 8'h75;
ROM_MEM[2880] = 8'h56;
ROM_MEM[2881] = 8'hEE;
ROM_MEM[2882] = 8'h58;
ROM_MEM[2883] = 8'h89;
ROM_MEM[2884] = 8'h32;
ROM_MEM[2885] = 8'h96;
ROM_MEM[2886] = 8'h1E;
ROM_MEM[2887] = 8'h78;
ROM_MEM[2888] = 8'hA3;
ROM_MEM[2889] = 8'h38;
ROM_MEM[2890] = 8'hF1;
ROM_MEM[2891] = 8'h5A;
ROM_MEM[2892] = 8'h7A;
ROM_MEM[2893] = 8'h94;
ROM_MEM[2894] = 8'hF5;
ROM_MEM[2895] = 8'h91;
ROM_MEM[2896] = 8'hC6;
ROM_MEM[2897] = 8'h63;
ROM_MEM[2898] = 8'h69;
ROM_MEM[2899] = 8'h81;
ROM_MEM[2900] = 8'hD7;
ROM_MEM[2901] = 8'hCB;
ROM_MEM[2902] = 8'h12;
ROM_MEM[2903] = 8'hB7;
ROM_MEM[2904] = 8'hA5;
ROM_MEM[2905] = 8'h79;
ROM_MEM[2906] = 8'hDE;
ROM_MEM[2907] = 8'h68;
ROM_MEM[2908] = 8'h75;
ROM_MEM[2909] = 8'hD8;
ROM_MEM[2910] = 8'hE6;
ROM_MEM[2911] = 8'h9E;
ROM_MEM[2912] = 8'h79;
ROM_MEM[2913] = 8'h3C;
ROM_MEM[2914] = 8'hC3;
ROM_MEM[2915] = 8'h66;
ROM_MEM[2916] = 8'h9B;
ROM_MEM[2917] = 8'h47;
ROM_MEM[2918] = 8'hD5;
ROM_MEM[2919] = 8'h92;
ROM_MEM[2920] = 8'hCC;
ROM_MEM[2921] = 8'h98;
ROM_MEM[2922] = 8'h6D;
ROM_MEM[2923] = 8'hE9;
ROM_MEM[2924] = 8'hC3;
ROM_MEM[2925] = 8'h12;
ROM_MEM[2926] = 8'h23;
ROM_MEM[2927] = 8'h13;
ROM_MEM[2928] = 8'h95;
ROM_MEM[2929] = 8'hB5;
ROM_MEM[2930] = 8'h57;
ROM_MEM[2931] = 8'h09;
ROM_MEM[2932] = 8'hCC;
ROM_MEM[2933] = 8'hAA;
ROM_MEM[2934] = 8'h55;
ROM_MEM[2935] = 8'hB6;
ROM_MEM[2936] = 8'h5E;
ROM_MEM[2937] = 8'hD8;
ROM_MEM[2938] = 8'hA5;
ROM_MEM[2939] = 8'h2B;
ROM_MEM[2940] = 8'h46;
ROM_MEM[2941] = 8'hDB;
ROM_MEM[2942] = 8'h5B;
ROM_MEM[2943] = 8'hA0;
ROM_MEM[2944] = 8'hF4;
ROM_MEM[2945] = 8'h4E;
ROM_MEM[2946] = 8'h53;
ROM_MEM[2947] = 8'h6C;
ROM_MEM[2948] = 8'h6F;
ROM_MEM[2949] = 8'h59;
ROM_MEM[2950] = 8'h5C;
ROM_MEM[2951] = 8'h3A;
ROM_MEM[2952] = 8'h2D;
ROM_MEM[2953] = 8'h9A;
ROM_MEM[2954] = 8'hAD;
ROM_MEM[2955] = 8'h16;
ROM_MEM[2956] = 8'h6E;
ROM_MEM[2957] = 8'hDD;
ROM_MEM[2958] = 8'hB2;
ROM_MEM[2959] = 8'h78;
ROM_MEM[2960] = 8'h96;
ROM_MEM[2961] = 8'h56;
ROM_MEM[2962] = 8'h35;
ROM_MEM[2963] = 8'hB5;
ROM_MEM[2964] = 8'hB3;
ROM_MEM[2965] = 8'hE1;
ROM_MEM[2966] = 8'h19;
ROM_MEM[2967] = 8'h5A;
ROM_MEM[2968] = 8'hD1;
ROM_MEM[2969] = 8'h92;
ROM_MEM[2970] = 8'h8D;
ROM_MEM[2971] = 8'h5A;
ROM_MEM[2972] = 8'hA7;
ROM_MEM[2973] = 8'hEB;
ROM_MEM[2974] = 8'h45;
ROM_MEM[2975] = 8'h53;
ROM_MEM[2976] = 8'hC6;
ROM_MEM[2977] = 8'h66;
ROM_MEM[2978] = 8'h9D;
ROM_MEM[2979] = 8'hBE;
ROM_MEM[2980] = 8'h57;
ROM_MEM[2981] = 8'h09;
ROM_MEM[2982] = 8'h19;
ROM_MEM[2983] = 8'h59;
ROM_MEM[2984] = 8'h3C;
ROM_MEM[2985] = 8'h86;
ROM_MEM[2986] = 8'h16;
ROM_MEM[2987] = 8'hB9;
ROM_MEM[2988] = 8'hB4;
ROM_MEM[2989] = 8'h25;
ROM_MEM[2990] = 8'h62;
ROM_MEM[2991] = 8'h1B;
ROM_MEM[2992] = 8'h5B;
ROM_MEM[2993] = 8'hA2;
ROM_MEM[2994] = 8'hE4;
ROM_MEM[2995] = 8'hF0;
ROM_MEM[2996] = 8'h88;
ROM_MEM[2997] = 8'h6D;
ROM_MEM[2998] = 8'hEC;
ROM_MEM[2999] = 8'h91;
ROM_MEM[3000] = 8'h42;
ROM_MEM[3001] = 8'h3C;
ROM_MEM[3002] = 8'h22;
ROM_MEM[3003] = 8'hB5;
ROM_MEM[3004] = 8'h7E;
ROM_MEM[3005] = 8'h04;
ROM_MEM[3006] = 8'h74;
ROM_MEM[3007] = 8'h1C;
ROM_MEM[3008] = 8'hAF;
ROM_MEM[3009] = 8'hDC;
ROM_MEM[3010] = 8'hFA;
ROM_MEM[3011] = 8'h11;
ROM_MEM[3012] = 8'hC8;
ROM_MEM[3013] = 8'h60;
ROM_MEM[3014] = 8'hFC;
ROM_MEM[3015] = 8'h76;
ROM_MEM[3016] = 8'hEB;
ROM_MEM[3017] = 8'h9A;
ROM_MEM[3018] = 8'h23;
ROM_MEM[3019] = 8'h85;
ROM_MEM[3020] = 8'h8B;
ROM_MEM[3021] = 8'hC6;
ROM_MEM[3022] = 8'hA5;
ROM_MEM[3023] = 8'h4D;
ROM_MEM[3024] = 8'h86;
ROM_MEM[3025] = 8'hDC;
ROM_MEM[3026] = 8'h57;
ROM_MEM[3027] = 8'h92;
ROM_MEM[3028] = 8'h94;
ROM_MEM[3029] = 8'h36;
ROM_MEM[3030] = 8'h09;
ROM_MEM[3031] = 8'h2E;
ROM_MEM[3032] = 8'h5B;
ROM_MEM[3033] = 8'h71;
ROM_MEM[3034] = 8'h53;
ROM_MEM[3035] = 8'hBA;
ROM_MEM[3036] = 8'hA0;
ROM_MEM[3037] = 8'h78;
ROM_MEM[3038] = 8'hA2;
ROM_MEM[3039] = 8'hC5;
ROM_MEM[3040] = 8'h6B;
ROM_MEM[3041] = 8'hE9;
ROM_MEM[3042] = 8'hB2;
ROM_MEM[3043] = 8'h82;
ROM_MEM[3044] = 8'h0E;
ROM_MEM[3045] = 8'h0B;
ROM_MEM[3046] = 8'h37;
ROM_MEM[3047] = 8'hA1;
ROM_MEM[3048] = 8'hAF;
ROM_MEM[3049] = 8'h1A;
ROM_MEM[3050] = 8'hAA;
ROM_MEM[3051] = 8'h2A;
ROM_MEM[3052] = 8'h6C;
ROM_MEM[3053] = 8'h8F;
ROM_MEM[3054] = 8'hBE;
ROM_MEM[3055] = 8'h05;
ROM_MEM[3056] = 8'h70;
ROM_MEM[3057] = 8'hCA;
ROM_MEM[3058] = 8'h48;
ROM_MEM[3059] = 8'h74;
ROM_MEM[3060] = 8'hC6;
ROM_MEM[3061] = 8'hDE;
ROM_MEM[3062] = 8'hA8;
ROM_MEM[3063] = 8'hA4;
ROM_MEM[3064] = 8'hD5;
ROM_MEM[3065] = 8'hD4;
ROM_MEM[3066] = 8'h5A;
ROM_MEM[3067] = 8'hAA;
ROM_MEM[3068] = 8'hE7;
ROM_MEM[3069] = 8'hB5;
ROM_MEM[3070] = 8'hD1;
ROM_MEM[3071] = 8'h50;
ROM_MEM[3072] = 8'h63;
ROM_MEM[3073] = 8'hAB;
ROM_MEM[3074] = 8'h41;
ROM_MEM[3075] = 8'h47;
ROM_MEM[3076] = 8'h4B;
ROM_MEM[3077] = 8'h2B;
ROM_MEM[3078] = 8'hB7;
ROM_MEM[3079] = 8'hA3;
ROM_MEM[3080] = 8'h38;
ROM_MEM[3081] = 8'hBD;
ROM_MEM[3082] = 8'h1C;
ROM_MEM[3083] = 8'hAA;
ROM_MEM[3084] = 8'hD4;
ROM_MEM[3085] = 8'hCE;
ROM_MEM[3086] = 8'hE2;
ROM_MEM[3087] = 8'h7D;
ROM_MEM[3088] = 8'hBD;
ROM_MEM[3089] = 8'hB9;
ROM_MEM[3090] = 8'hF1;
ROM_MEM[3091] = 8'hB8;
ROM_MEM[3092] = 8'h9A;
ROM_MEM[3093] = 8'h93;
ROM_MEM[3094] = 8'h89;
ROM_MEM[3095] = 8'hA5;
ROM_MEM[3096] = 8'hD8;
ROM_MEM[3097] = 8'hED;
ROM_MEM[3098] = 8'hCA;
ROM_MEM[3099] = 8'h36;
ROM_MEM[3100] = 8'h2E;
ROM_MEM[3101] = 8'h12;
ROM_MEM[3102] = 8'h13;
ROM_MEM[3103] = 8'h97;
ROM_MEM[3104] = 8'hAB;
ROM_MEM[3105] = 8'h1A;
ROM_MEM[3106] = 8'hDB;
ROM_MEM[3107] = 8'h1C;
ROM_MEM[3108] = 8'h64;
ROM_MEM[3109] = 8'h5D;
ROM_MEM[3110] = 8'hEE;
ROM_MEM[3111] = 8'hE1;
ROM_MEM[3112] = 8'hA8;
ROM_MEM[3113] = 8'hE2;
ROM_MEM[3114] = 8'h50;
ROM_MEM[3115] = 8'h6D;
ROM_MEM[3116] = 8'hB8;
ROM_MEM[3117] = 8'hBB;
ROM_MEM[3118] = 8'hA4;
ROM_MEM[3119] = 8'h8B;
ROM_MEM[3120] = 8'h14;
ROM_MEM[3121] = 8'h35;
ROM_MEM[3122] = 8'hE9;
ROM_MEM[3123] = 8'hCE;
ROM_MEM[3124] = 8'hDC;
ROM_MEM[3125] = 8'hD6;
ROM_MEM[3126] = 8'h45;
ROM_MEM[3127] = 8'hD5;
ROM_MEM[3128] = 8'hA6;
ROM_MEM[3129] = 8'hBB;
ROM_MEM[3130] = 8'h72;
ROM_MEM[3131] = 8'hDE;
ROM_MEM[3132] = 8'h36;
ROM_MEM[3133] = 8'h51;
ROM_MEM[3134] = 8'h14;
ROM_MEM[3135] = 8'hEE;
ROM_MEM[3136] = 8'hC2;
ROM_MEM[3137] = 8'hF9;
ROM_MEM[3138] = 8'h4A;
ROM_MEM[3139] = 8'hD5;
ROM_MEM[3140] = 8'h91;
ROM_MEM[3141] = 8'hBD;
ROM_MEM[3142] = 8'h1F;
ROM_MEM[3143] = 8'hE0;
ROM_MEM[3144] = 8'hF5;
ROM_MEM[3145] = 8'hB2;
ROM_MEM[3146] = 8'hAE;
ROM_MEM[3147] = 8'h8F;
ROM_MEM[3148] = 8'hD4;
ROM_MEM[3149] = 8'h47;
ROM_MEM[3150] = 8'hCD;
ROM_MEM[3151] = 8'h9C;
ROM_MEM[3152] = 8'h26;
ROM_MEM[3153] = 8'h4B;
ROM_MEM[3154] = 8'hC6;
ROM_MEM[3155] = 8'h49;
ROM_MEM[3156] = 8'h8A;
ROM_MEM[3157] = 8'h4E;
ROM_MEM[3158] = 8'hDD;
ROM_MEM[3159] = 8'hD4;
ROM_MEM[3160] = 8'h60;
ROM_MEM[3161] = 8'hA7;
ROM_MEM[3162] = 8'h28;
ROM_MEM[3163] = 8'hDA;
ROM_MEM[3164] = 8'hF1;
ROM_MEM[3165] = 8'h50;
ROM_MEM[3166] = 8'h82;
ROM_MEM[3167] = 8'hED;
ROM_MEM[3168] = 8'hE0;
ROM_MEM[3169] = 8'hAC;
ROM_MEM[3170] = 8'h28;
ROM_MEM[3171] = 8'h46;
ROM_MEM[3172] = 8'h89;
ROM_MEM[3173] = 8'hAC;
ROM_MEM[3174] = 8'h2A;
ROM_MEM[3175] = 8'hDC;
ROM_MEM[3176] = 8'h12;
ROM_MEM[3177] = 8'h2B;
ROM_MEM[3178] = 8'h25;
ROM_MEM[3179] = 8'hD2;
ROM_MEM[3180] = 8'hAC;
ROM_MEM[3181] = 8'h50;
ROM_MEM[3182] = 8'hB7;
ROM_MEM[3183] = 8'h6D;
ROM_MEM[3184] = 8'h80;
ROM_MEM[3185] = 8'h52;
ROM_MEM[3186] = 8'h58;
ROM_MEM[3187] = 8'h87;
ROM_MEM[3188] = 8'hDE;
ROM_MEM[3189] = 8'h56;
ROM_MEM[3190] = 8'h08;
ROM_MEM[3191] = 8'h6B;
ROM_MEM[3192] = 8'h38;
ROM_MEM[3193] = 8'h39;
ROM_MEM[3194] = 8'h5E;
ROM_MEM[3195] = 8'h11;
ROM_MEM[3196] = 8'hE2;
ROM_MEM[3197] = 8'hE9;
ROM_MEM[3198] = 8'h45;
ROM_MEM[3199] = 8'hB9;
ROM_MEM[3200] = 8'h04;
ROM_MEM[3201] = 8'h89;
ROM_MEM[3202] = 8'hB0;
ROM_MEM[3203] = 8'h59;
ROM_MEM[3204] = 8'h94;
ROM_MEM[3205] = 8'h15;
ROM_MEM[3206] = 8'h30;
ROM_MEM[3207] = 8'h7E;
ROM_MEM[3208] = 8'hA2;
ROM_MEM[3209] = 8'hA2;
ROM_MEM[3210] = 8'h9E;
ROM_MEM[3211] = 8'h25;
ROM_MEM[3212] = 8'h35;
ROM_MEM[3213] = 8'h05;
ROM_MEM[3214] = 8'hCD;
ROM_MEM[3215] = 8'h2B;
ROM_MEM[3216] = 8'h8B;
ROM_MEM[3217] = 8'h46;
ROM_MEM[3218] = 8'h9C;
ROM_MEM[3219] = 8'hE1;
ROM_MEM[3220] = 8'h27;
ROM_MEM[3221] = 8'h2D;
ROM_MEM[3222] = 8'hAE;
ROM_MEM[3223] = 8'h35;
ROM_MEM[3224] = 8'h32;
ROM_MEM[3225] = 8'h4F;
ROM_MEM[3226] = 8'h50;
ROM_MEM[3227] = 8'h94;
ROM_MEM[3228] = 8'h84;
ROM_MEM[3229] = 8'hD6;
ROM_MEM[3230] = 8'h28;
ROM_MEM[3231] = 8'h5C;
ROM_MEM[3232] = 8'h61;
ROM_MEM[3233] = 8'hA6;
ROM_MEM[3234] = 8'hEA;
ROM_MEM[3235] = 8'hA9;
ROM_MEM[3236] = 8'h2D;
ROM_MEM[3237] = 8'h69;
ROM_MEM[3238] = 8'h45;
ROM_MEM[3239] = 8'h83;
ROM_MEM[3240] = 8'h1B;
ROM_MEM[3241] = 8'hB3;
ROM_MEM[3242] = 8'h44;
ROM_MEM[3243] = 8'h92;
ROM_MEM[3244] = 8'h11;
ROM_MEM[3245] = 8'h2E;
ROM_MEM[3246] = 8'h65;
ROM_MEM[3247] = 8'h2C;
ROM_MEM[3248] = 8'h92;
ROM_MEM[3249] = 8'h89;
ROM_MEM[3250] = 8'h47;
ROM_MEM[3251] = 8'hB8;
ROM_MEM[3252] = 8'hDC;
ROM_MEM[3253] = 8'hB8;
ROM_MEM[3254] = 8'h91;
ROM_MEM[3255] = 8'hD8;
ROM_MEM[3256] = 8'h0E;
ROM_MEM[3257] = 8'hC0;
ROM_MEM[3258] = 8'h14;
ROM_MEM[3259] = 8'hCC;
ROM_MEM[3260] = 8'h01;
ROM_MEM[3261] = 8'h98;
ROM_MEM[3262] = 8'h9C;
ROM_MEM[3263] = 8'h38;
ROM_MEM[3264] = 8'h01;
ROM_MEM[3265] = 8'h47;
ROM_MEM[3266] = 8'h39;
ROM_MEM[3267] = 8'h15;
ROM_MEM[3268] = 8'h60;
ROM_MEM[3269] = 8'h48;
ROM_MEM[3270] = 8'h93;
ROM_MEM[3271] = 8'hA5;
ROM_MEM[3272] = 8'h54;
ROM_MEM[3273] = 8'h65;
ROM_MEM[3274] = 8'hAE;
ROM_MEM[3275] = 8'h9E;
ROM_MEM[3276] = 8'h8A;
ROM_MEM[3277] = 8'h8F;
ROM_MEM[3278] = 8'h9C;
ROM_MEM[3279] = 8'h6C;
ROM_MEM[3280] = 8'hBA;
ROM_MEM[3281] = 8'h66;
ROM_MEM[3282] = 8'h2A;
ROM_MEM[3283] = 8'h3A;
ROM_MEM[3284] = 8'h72;
ROM_MEM[3285] = 8'h36;
ROM_MEM[3286] = 8'h5E;
ROM_MEM[3287] = 8'hE2;
ROM_MEM[3288] = 8'h66;
ROM_MEM[3289] = 8'hF3;
ROM_MEM[3290] = 8'h88;
ROM_MEM[3291] = 8'hD5;
ROM_MEM[3292] = 8'hC5;
ROM_MEM[3293] = 8'h48;
ROM_MEM[3294] = 8'h9A;
ROM_MEM[3295] = 8'hED;
ROM_MEM[3296] = 8'h23;
ROM_MEM[3297] = 8'h34;
ROM_MEM[3298] = 8'h17;
ROM_MEM[3299] = 8'h4D;
ROM_MEM[3300] = 8'h29;
ROM_MEM[3301] = 8'hB2;
ROM_MEM[3302] = 8'h0F;
ROM_MEM[3303] = 8'hDB;
ROM_MEM[3304] = 8'h9D;
ROM_MEM[3305] = 8'h17;
ROM_MEM[3306] = 8'hA7;
ROM_MEM[3307] = 8'h3B;
ROM_MEM[3308] = 8'h39;
ROM_MEM[3309] = 8'h74;
ROM_MEM[3310] = 8'hF7;
ROM_MEM[3311] = 8'h11;
ROM_MEM[3312] = 8'h34;
ROM_MEM[3313] = 8'h1E;
ROM_MEM[3314] = 8'hFB;
ROM_MEM[3315] = 8'hD0;
ROM_MEM[3316] = 8'hAD;
ROM_MEM[3317] = 8'h9A;
ROM_MEM[3318] = 8'h4B;
ROM_MEM[3319] = 8'h77;
ROM_MEM[3320] = 8'hEC;
ROM_MEM[3321] = 8'h43;
ROM_MEM[3322] = 8'hF7;
ROM_MEM[3323] = 8'h64;
ROM_MEM[3324] = 8'h26;
ROM_MEM[3325] = 8'hD9;
ROM_MEM[3326] = 8'hAD;
ROM_MEM[3327] = 8'h0E;
ROM_MEM[3328] = 8'hDB;
ROM_MEM[3329] = 8'hAD;
ROM_MEM[3330] = 8'h98;
ROM_MEM[3331] = 8'h5D;
ROM_MEM[3332] = 8'hC7;
ROM_MEM[3333] = 8'h3A;
ROM_MEM[3334] = 8'hC2;
ROM_MEM[3335] = 8'h70;
ROM_MEM[3336] = 8'hA2;
ROM_MEM[3337] = 8'hD8;
ROM_MEM[3338] = 8'h69;
ROM_MEM[3339] = 8'h6B;
ROM_MEM[3340] = 8'h98;
ROM_MEM[3341] = 8'h8B;
ROM_MEM[3342] = 8'h27;
ROM_MEM[3343] = 8'hB3;
ROM_MEM[3344] = 8'h55;
ROM_MEM[3345] = 8'hAD;
ROM_MEM[3346] = 8'hE5;
ROM_MEM[3347] = 8'h6F;
ROM_MEM[3348] = 8'h6E;
ROM_MEM[3349] = 8'h4C;
ROM_MEM[3350] = 8'h14;
ROM_MEM[3351] = 8'h89;
ROM_MEM[3352] = 8'h57;
ROM_MEM[3353] = 8'hB4;
ROM_MEM[3354] = 8'hA8;
ROM_MEM[3355] = 8'hB2;
ROM_MEM[3356] = 8'h4A;
ROM_MEM[3357] = 8'hC4;
ROM_MEM[3358] = 8'h3E;
ROM_MEM[3359] = 8'h41;
ROM_MEM[3360] = 8'h57;
ROM_MEM[3361] = 8'h62;
ROM_MEM[3362] = 8'hCA;
ROM_MEM[3363] = 8'hE9;
ROM_MEM[3364] = 8'hE8;
ROM_MEM[3365] = 8'h44;
ROM_MEM[3366] = 8'h4D;
ROM_MEM[3367] = 8'h71;
ROM_MEM[3368] = 8'h72;
ROM_MEM[3369] = 8'h96;
ROM_MEM[3370] = 8'hCD;
ROM_MEM[3371] = 8'h15;
ROM_MEM[3372] = 8'h67;
ROM_MEM[3373] = 8'hA1;
ROM_MEM[3374] = 8'h49;
ROM_MEM[3375] = 8'hDE;
ROM_MEM[3376] = 8'hB6;
ROM_MEM[3377] = 8'h18;
ROM_MEM[3378] = 8'hC0;
ROM_MEM[3379] = 8'hB4;
ROM_MEM[3380] = 8'h97;
ROM_MEM[3381] = 8'h02;
ROM_MEM[3382] = 8'hA8;
ROM_MEM[3383] = 8'h8D;
ROM_MEM[3384] = 8'h38;
ROM_MEM[3385] = 8'h69;
ROM_MEM[3386] = 8'hF5;
ROM_MEM[3387] = 8'h6A;
ROM_MEM[3388] = 8'hD4;
ROM_MEM[3389] = 8'hED;
ROM_MEM[3390] = 8'hF0;
ROM_MEM[3391] = 8'hE4;
ROM_MEM[3392] = 8'hCD;
ROM_MEM[3393] = 8'h49;
ROM_MEM[3394] = 8'hE8;
ROM_MEM[3395] = 8'hB4;
ROM_MEM[3396] = 8'hCD;
ROM_MEM[3397] = 8'h53;
ROM_MEM[3398] = 8'h94;
ROM_MEM[3399] = 8'hC2;
ROM_MEM[3400] = 8'h1E;
ROM_MEM[3401] = 8'h5B;
ROM_MEM[3402] = 8'hB2;
ROM_MEM[3403] = 8'h4E;
ROM_MEM[3404] = 8'hDE;
ROM_MEM[3405] = 8'hAA;
ROM_MEM[3406] = 8'h89;
ROM_MEM[3407] = 8'h56;
ROM_MEM[3408] = 8'h39;
ROM_MEM[3409] = 8'h3C;
ROM_MEM[3410] = 8'h65;
ROM_MEM[3411] = 8'hB1;
ROM_MEM[3412] = 8'h16;
ROM_MEM[3413] = 8'h91;
ROM_MEM[3414] = 8'h63;
ROM_MEM[3415] = 8'h25;
ROM_MEM[3416] = 8'hE4;
ROM_MEM[3417] = 8'h55;
ROM_MEM[3418] = 8'h9B;
ROM_MEM[3419] = 8'h59;
ROM_MEM[3420] = 8'h84;
ROM_MEM[3421] = 8'h68;
ROM_MEM[3422] = 8'h06;
ROM_MEM[3423] = 8'h48;
ROM_MEM[3424] = 8'hE5;
ROM_MEM[3425] = 8'h49;
ROM_MEM[3426] = 8'h00;
ROM_MEM[3427] = 8'h29;
ROM_MEM[3428] = 8'h23;
ROM_MEM[3429] = 8'h10;
ROM_MEM[3430] = 8'h20;
ROM_MEM[3431] = 8'h71;
ROM_MEM[3432] = 8'h98;
ROM_MEM[3433] = 8'h00;
ROM_MEM[3434] = 8'h0A;
ROM_MEM[3435] = 8'h67;
ROM_MEM[3436] = 8'h31;
ROM_MEM[3437] = 8'h40;
ROM_MEM[3438] = 8'h31;
ROM_MEM[3439] = 8'h6A;
ROM_MEM[3440] = 8'h2B;
ROM_MEM[3441] = 8'h6C;
ROM_MEM[3442] = 8'h41;
ROM_MEM[3443] = 8'h8D;
ROM_MEM[3444] = 8'h74;
ROM_MEM[3445] = 8'h1D;
ROM_MEM[3446] = 8'h9E;
ROM_MEM[3447] = 8'hA8;
ROM_MEM[3448] = 8'h79;
ROM_MEM[3449] = 8'h33;
ROM_MEM[3450] = 8'hF6;
ROM_MEM[3451] = 8'h8D;
ROM_MEM[3452] = 8'h79;
ROM_MEM[3453] = 8'hE2;
ROM_MEM[3454] = 8'h16;
ROM_MEM[3455] = 8'hD4;
ROM_MEM[3456] = 8'hA4;
ROM_MEM[3457] = 8'h26;
ROM_MEM[3458] = 8'hE1;
ROM_MEM[3459] = 8'h49;
ROM_MEM[3460] = 8'h7B;
ROM_MEM[3461] = 8'h31;
ROM_MEM[3462] = 8'hC3;
ROM_MEM[3463] = 8'hEA;
ROM_MEM[3464] = 8'h58;
ROM_MEM[3465] = 8'h27;
ROM_MEM[3466] = 8'hEB;
ROM_MEM[3467] = 8'h49;
ROM_MEM[3468] = 8'h0D;
ROM_MEM[3469] = 8'hBB;
ROM_MEM[3470] = 8'h6C;
ROM_MEM[3471] = 8'hAD;
ROM_MEM[3472] = 8'hBC;
ROM_MEM[3473] = 8'h27;
ROM_MEM[3474] = 8'h16;
ROM_MEM[3475] = 8'hAD;
ROM_MEM[3476] = 8'h92;
ROM_MEM[3477] = 8'h38;
ROM_MEM[3478] = 8'hCA;
ROM_MEM[3479] = 8'h11;
ROM_MEM[3480] = 8'h48;
ROM_MEM[3481] = 8'h3D;
ROM_MEM[3482] = 8'h43;
ROM_MEM[3483] = 8'h52;
ROM_MEM[3484] = 8'hAA;
ROM_MEM[3485] = 8'h9A;
ROM_MEM[3486] = 8'h41;
ROM_MEM[3487] = 8'hF7;
ROM_MEM[3488] = 8'h72;
ROM_MEM[3489] = 8'h8B;
ROM_MEM[3490] = 8'hA1;
ROM_MEM[3491] = 8'hA9;
ROM_MEM[3492] = 8'h9A;
ROM_MEM[3493] = 8'hCC;
ROM_MEM[3494] = 8'hD2;
ROM_MEM[3495] = 8'h93;
ROM_MEM[3496] = 8'h30;
ROM_MEM[3497] = 8'h40;
ROM_MEM[3498] = 8'h48;
ROM_MEM[3499] = 8'h1B;
ROM_MEM[3500] = 8'hD7;
ROM_MEM[3501] = 8'h75;
ROM_MEM[3502] = 8'h23;
ROM_MEM[3503] = 8'h2A;
ROM_MEM[3504] = 8'hE6;
ROM_MEM[3505] = 8'h76;
ROM_MEM[3506] = 8'h08;
ROM_MEM[3507] = 8'hC0;
ROM_MEM[3508] = 8'h65;
ROM_MEM[3509] = 8'hD4;
ROM_MEM[3510] = 8'h03;
ROM_MEM[3511] = 8'h86;
ROM_MEM[3512] = 8'h34;
ROM_MEM[3513] = 8'h29;
ROM_MEM[3514] = 8'h04;
ROM_MEM[3515] = 8'h88;
ROM_MEM[3516] = 8'h98;
ROM_MEM[3517] = 8'h84;
ROM_MEM[3518] = 8'h00;
ROM_MEM[3519] = 8'h99;
ROM_MEM[3520] = 8'h20;
ROM_MEM[3521] = 8'h11;
ROM_MEM[3522] = 8'hA0;
ROM_MEM[3523] = 8'h71;
ROM_MEM[3524] = 8'h62;
ROM_MEM[3525] = 8'h06;
ROM_MEM[3526] = 8'h34;
ROM_MEM[3527] = 8'hC1;
ROM_MEM[3528] = 8'hCC;
ROM_MEM[3529] = 8'h80;
ROM_MEM[3530] = 8'h2E;
ROM_MEM[3531] = 8'h58;
ROM_MEM[3532] = 8'h10;
ROM_MEM[3533] = 8'h90;
ROM_MEM[3534] = 8'h18;
ROM_MEM[3535] = 8'h09;
ROM_MEM[3536] = 8'h02;
ROM_MEM[3537] = 8'h3C;
ROM_MEM[3538] = 8'h52;
ROM_MEM[3539] = 8'h23;
ROM_MEM[3540] = 8'h80;
ROM_MEM[3541] = 8'hE5;
ROM_MEM[3542] = 8'h1E;
ROM_MEM[3543] = 8'hAD;
ROM_MEM[3544] = 8'h6D;
ROM_MEM[3545] = 8'h45;
ROM_MEM[3546] = 8'h8D;
ROM_MEM[3547] = 8'h3C;
ROM_MEM[3548] = 8'h3B;
ROM_MEM[3549] = 8'hAD;
ROM_MEM[3550] = 8'hB6;
ROM_MEM[3551] = 8'h4D;
ROM_MEM[3552] = 8'h6F;
ROM_MEM[3553] = 8'h10;
ROM_MEM[3554] = 8'h5A;
ROM_MEM[3555] = 8'hB3;
ROM_MEM[3556] = 8'hDA;
ROM_MEM[3557] = 8'h36;
ROM_MEM[3558] = 8'h39;
ROM_MEM[3559] = 8'hA1;
ROM_MEM[3560] = 8'hE2;
ROM_MEM[3561] = 8'hCD;
ROM_MEM[3562] = 8'hA9;
ROM_MEM[3563] = 8'hDB;
ROM_MEM[3564] = 8'hE0;
ROM_MEM[3565] = 8'h84;
ROM_MEM[3566] = 8'hCE;
ROM_MEM[3567] = 8'h35;
ROM_MEM[3568] = 8'hA3;
ROM_MEM[3569] = 8'h6A;
ROM_MEM[3570] = 8'h8D;
ROM_MEM[3571] = 8'h02;
ROM_MEM[3572] = 8'h27;
ROM_MEM[3573] = 8'hBF;
ROM_MEM[3574] = 8'hAC;
ROM_MEM[3575] = 8'hBC;
ROM_MEM[3576] = 8'h0F;
ROM_MEM[3577] = 8'h0A;
ROM_MEM[3578] = 8'h98;
ROM_MEM[3579] = 8'h5C;
ROM_MEM[3580] = 8'hB5;
ROM_MEM[3581] = 8'hF2;
ROM_MEM[3582] = 8'h7E;
ROM_MEM[3583] = 8'h34;
ROM_MEM[3584] = 8'h21;
ROM_MEM[3585] = 8'h64;
ROM_MEM[3586] = 8'hF5;
ROM_MEM[3587] = 8'h4A;
ROM_MEM[3588] = 8'h7B;
ROM_MEM[3589] = 8'h45;
ROM_MEM[3590] = 8'hC7;
ROM_MEM[3591] = 8'hAB;
ROM_MEM[3592] = 8'h4D;
ROM_MEM[3593] = 8'h2B;
ROM_MEM[3594] = 8'hE9;
ROM_MEM[3595] = 8'h0D;
ROM_MEM[3596] = 8'h1D;
ROM_MEM[3597] = 8'h37;
ROM_MEM[3598] = 8'h37;
ROM_MEM[3599] = 8'h8E;
ROM_MEM[3600] = 8'hB8;
ROM_MEM[3601] = 8'h77;
ROM_MEM[3602] = 8'h74;
ROM_MEM[3603] = 8'hDC;
ROM_MEM[3604] = 8'h5C;
ROM_MEM[3605] = 8'h58;
ROM_MEM[3606] = 8'hE2;
ROM_MEM[3607] = 8'h56;
ROM_MEM[3608] = 8'h20;
ROM_MEM[3609] = 8'h65;
ROM_MEM[3610] = 8'hBB;
ROM_MEM[3611] = 8'h51;
ROM_MEM[3612] = 8'h49;
ROM_MEM[3613] = 8'h9A;
ROM_MEM[3614] = 8'h87;
ROM_MEM[3615] = 8'hB4;
ROM_MEM[3616] = 8'hAB;
ROM_MEM[3617] = 8'h96;
ROM_MEM[3618] = 8'hAD;
ROM_MEM[3619] = 8'hEF;
ROM_MEM[3620] = 8'h9D;
ROM_MEM[3621] = 8'h03;
ROM_MEM[3622] = 8'hCA;
ROM_MEM[3623] = 8'h17;
ROM_MEM[3624] = 8'h8D;
ROM_MEM[3625] = 8'hBE;
ROM_MEM[3626] = 8'h0F;
ROM_MEM[3627] = 8'h4D;
ROM_MEM[3628] = 8'h28;
ROM_MEM[3629] = 8'hBB;
ROM_MEM[3630] = 8'h35;
ROM_MEM[3631] = 8'hFA;
ROM_MEM[3632] = 8'h36;
ROM_MEM[3633] = 8'h35;
ROM_MEM[3634] = 8'hA1;
ROM_MEM[3635] = 8'h7C;
ROM_MEM[3636] = 8'h56;
ROM_MEM[3637] = 8'h19;
ROM_MEM[3638] = 8'h4A;
ROM_MEM[3639] = 8'h00;
ROM_MEM[3640] = 8'h97;
ROM_MEM[3641] = 8'h2E;
ROM_MEM[3642] = 8'hDB;
ROM_MEM[3643] = 8'hA5;
ROM_MEM[3644] = 8'hAF;
ROM_MEM[3645] = 8'h11;
ROM_MEM[3646] = 8'h92;
ROM_MEM[3647] = 8'hB3;
ROM_MEM[3648] = 8'h12;
ROM_MEM[3649] = 8'hAF;
ROM_MEM[3650] = 8'hBE;
ROM_MEM[3651] = 8'h15;
ROM_MEM[3652] = 8'h2A;
ROM_MEM[3653] = 8'h6C;
ROM_MEM[3654] = 8'hAF;
ROM_MEM[3655] = 8'hBD;
ROM_MEM[3656] = 8'hC6;
ROM_MEM[3657] = 8'hDE;
ROM_MEM[3658] = 8'hA9;
ROM_MEM[3659] = 8'hB1;
ROM_MEM[3660] = 8'hBC;
ROM_MEM[3661] = 8'h4D;
ROM_MEM[3662] = 8'h0A;
ROM_MEM[3663] = 8'hAB;
ROM_MEM[3664] = 8'hC7;
ROM_MEM[3665] = 8'hD6;
ROM_MEM[3666] = 8'hEA;
ROM_MEM[3667] = 8'hC6;
ROM_MEM[3668] = 8'h61;
ROM_MEM[3669] = 8'h2C;
ROM_MEM[3670] = 8'h0E;
ROM_MEM[3671] = 8'h3D;
ROM_MEM[3672] = 8'hAC;
ROM_MEM[3673] = 8'h22;
ROM_MEM[3674] = 8'h11;
ROM_MEM[3675] = 8'hC0;
ROM_MEM[3676] = 8'h18;
ROM_MEM[3677] = 8'h4B;
ROM_MEM[3678] = 8'h02;
ROM_MEM[3679] = 8'h68;
ROM_MEM[3680] = 8'hED;
ROM_MEM[3681] = 8'h61;
ROM_MEM[3682] = 8'h80;
ROM_MEM[3683] = 8'h64;
ROM_MEM[3684] = 8'h28;
ROM_MEM[3685] = 8'h4A;
ROM_MEM[3686] = 8'h55;
ROM_MEM[3687] = 8'h02;
ROM_MEM[3688] = 8'h8F;
ROM_MEM[3689] = 8'h65;
ROM_MEM[3690] = 8'hC6;
ROM_MEM[3691] = 8'h3A;
ROM_MEM[3692] = 8'h65;
ROM_MEM[3693] = 8'h09;
ROM_MEM[3694] = 8'hDC;
ROM_MEM[3695] = 8'hBA;
ROM_MEM[3696] = 8'h16;
ROM_MEM[3697] = 8'hFB;
ROM_MEM[3698] = 8'h54;
ROM_MEM[3699] = 8'hAD;
ROM_MEM[3700] = 8'hF3;
ROM_MEM[3701] = 8'h48;
ROM_MEM[3702] = 8'h79;
ROM_MEM[3703] = 8'hEB;
ROM_MEM[3704] = 8'h93;
ROM_MEM[3705] = 8'hF7;
ROM_MEM[3706] = 8'hC5;
ROM_MEM[3707] = 8'hC5;
ROM_MEM[3708] = 8'hAD;
ROM_MEM[3709] = 8'h4D;
ROM_MEM[3710] = 8'h5A;
ROM_MEM[3711] = 8'h5E;
ROM_MEM[3712] = 8'h13;
ROM_MEM[3713] = 8'h15;
ROM_MEM[3714] = 8'h4F;
ROM_MEM[3715] = 8'h5A;
ROM_MEM[3716] = 8'h4A;
ROM_MEM[3717] = 8'h79;
ROM_MEM[3718] = 8'hCD;
ROM_MEM[3719] = 8'h92;
ROM_MEM[3720] = 8'h92;
ROM_MEM[3721] = 8'hE1;
ROM_MEM[3722] = 8'h98;
ROM_MEM[3723] = 8'h01;
ROM_MEM[3724] = 8'hD2;
ROM_MEM[3725] = 8'h49;
ROM_MEM[3726] = 8'h12;
ROM_MEM[3727] = 8'hC0;
ROM_MEM[3728] = 8'h2B;
ROM_MEM[3729] = 8'h0D;
ROM_MEM[3730] = 8'h02;
ROM_MEM[3731] = 8'h78;
ROM_MEM[3732] = 8'h65;
ROM_MEM[3733] = 8'h46;
ROM_MEM[3734] = 8'h80;
ROM_MEM[3735] = 8'h60;
ROM_MEM[3736] = 8'h5D;
ROM_MEM[3737] = 8'h05;
ROM_MEM[3738] = 8'h90;
ROM_MEM[3739] = 8'h22;
ROM_MEM[3740] = 8'hBB;
ROM_MEM[3741] = 8'h02;
ROM_MEM[3742] = 8'h8A;
ROM_MEM[3743] = 8'hA1;
ROM_MEM[3744] = 8'h10;
ROM_MEM[3745] = 8'h40;
ROM_MEM[3746] = 8'hD6;
ROM_MEM[3747] = 8'hEC;
ROM_MEM[3748] = 8'h0C;
ROM_MEM[3749] = 8'h48;
ROM_MEM[3750] = 8'h8A;
ROM_MEM[3751] = 8'h23;
ROM_MEM[3752] = 8'h44;
ROM_MEM[3753] = 8'hD1;
ROM_MEM[3754] = 8'h48;
ROM_MEM[3755] = 8'h56;
ROM_MEM[3756] = 8'h45;
ROM_MEM[3757] = 8'hAC;
ROM_MEM[3758] = 8'h90;
ROM_MEM[3759] = 8'hDB;
ROM_MEM[3760] = 8'hD0;
ROM_MEM[3761] = 8'h9D;
ROM_MEM[3762] = 8'h6E;
ROM_MEM[3763] = 8'hB6;
ROM_MEM[3764] = 8'h4B;
ROM_MEM[3765] = 8'h61;
ROM_MEM[3766] = 8'h42;
ROM_MEM[3767] = 8'hAD;
ROM_MEM[3768] = 8'h07;
ROM_MEM[3769] = 8'h65;
ROM_MEM[3770] = 8'h29;
ROM_MEM[3771] = 8'hB9;
ROM_MEM[3772] = 8'h49;
ROM_MEM[3773] = 8'h75;
ROM_MEM[3774] = 8'h11;
ROM_MEM[3775] = 8'hEC;
ROM_MEM[3776] = 8'hA5;
ROM_MEM[3777] = 8'hE5;
ROM_MEM[3778] = 8'hCE;
ROM_MEM[3779] = 8'hE5;
ROM_MEM[3780] = 8'h79;
ROM_MEM[3781] = 8'h72;
ROM_MEM[3782] = 8'hEA;
ROM_MEM[3783] = 8'hD2;
ROM_MEM[3784] = 8'h06;
ROM_MEM[3785] = 8'h2B;
ROM_MEM[3786] = 8'h93;
ROM_MEM[3787] = 8'hAE;
ROM_MEM[3788] = 8'h8E;
ROM_MEM[3789] = 8'h4B;
ROM_MEM[3790] = 8'h57;
ROM_MEM[3791] = 8'h02;
ROM_MEM[3792] = 8'hA6;
ROM_MEM[3793] = 8'h78;
ROM_MEM[3794] = 8'hD8;
ROM_MEM[3795] = 8'h1A;
ROM_MEM[3796] = 8'h43;
ROM_MEM[3797] = 8'h89;
ROM_MEM[3798] = 8'h14;
ROM_MEM[3799] = 8'h9C;
ROM_MEM[3800] = 8'h5A;
ROM_MEM[3801] = 8'h3B;
ROM_MEM[3802] = 8'h00;
ROM_MEM[3803] = 8'hC9;
ROM_MEM[3804] = 8'h42;
ROM_MEM[3805] = 8'hB5;
ROM_MEM[3806] = 8'hBE;
ROM_MEM[3807] = 8'h2D;
ROM_MEM[3808] = 8'h71;
ROM_MEM[3809] = 8'h68;
ROM_MEM[3810] = 8'h6F;
ROM_MEM[3811] = 8'h95;
ROM_MEM[3812] = 8'hB2;
ROM_MEM[3813] = 8'h5E;
ROM_MEM[3814] = 8'hC8;
ROM_MEM[3815] = 8'hA1;
ROM_MEM[3816] = 8'hB2;
ROM_MEM[3817] = 8'h55;
ROM_MEM[3818] = 8'hDA;
ROM_MEM[3819] = 8'h7B;
ROM_MEM[3820] = 8'h57;
ROM_MEM[3821] = 8'h07;
ROM_MEM[3822] = 8'h89;
ROM_MEM[3823] = 8'h34;
ROM_MEM[3824] = 8'h0E;
ROM_MEM[3825] = 8'h68;
ROM_MEM[3826] = 8'h09;
ROM_MEM[3827] = 8'hDD;
ROM_MEM[3828] = 8'h00;
ROM_MEM[3829] = 8'h2D;
ROM_MEM[3830] = 8'h90;
ROM_MEM[3831] = 8'h29;
ROM_MEM[3832] = 8'h20;
ROM_MEM[3833] = 8'h49;
ROM_MEM[3834] = 8'hAA;
ROM_MEM[3835] = 8'h50;
ROM_MEM[3836] = 8'h35;
ROM_MEM[3837] = 8'h0B;
ROM_MEM[3838] = 8'h61;
ROM_MEM[3839] = 8'h11;
ROM_MEM[3840] = 8'h8E;
ROM_MEM[3841] = 8'hDD;
ROM_MEM[3842] = 8'h5A;
ROM_MEM[3843] = 8'h14;
ROM_MEM[3844] = 8'h78;
ROM_MEM[3845] = 8'h46;
ROM_MEM[3846] = 8'h45;
ROM_MEM[3847] = 8'h0E;
ROM_MEM[3848] = 8'h6B;
ROM_MEM[3849] = 8'h16;
ROM_MEM[3850] = 8'hE8;
ROM_MEM[3851] = 8'h19;
ROM_MEM[3852] = 8'h15;
ROM_MEM[3853] = 8'hD9;
ROM_MEM[3854] = 8'h6D;
ROM_MEM[3855] = 8'h89;
ROM_MEM[3856] = 8'h51;
ROM_MEM[3857] = 8'hB5;
ROM_MEM[3858] = 8'hBB;
ROM_MEM[3859] = 8'hED;
ROM_MEM[3860] = 8'hB0;
ROM_MEM[3861] = 8'h65;
ROM_MEM[3862] = 8'hC6;
ROM_MEM[3863] = 8'h5E;
ROM_MEM[3864] = 8'h11;
ROM_MEM[3865] = 8'h8E;
ROM_MEM[3866] = 8'hDD;
ROM_MEM[3867] = 8'h5E;
ROM_MEM[3868] = 8'h98;
ROM_MEM[3869] = 8'h98;
ROM_MEM[3870] = 8'h47;
ROM_MEM[3871] = 8'hD8;
ROM_MEM[3872] = 8'h36;
ROM_MEM[3873] = 8'h7B;
ROM_MEM[3874] = 8'h26;
ROM_MEM[3875] = 8'hA2;
ROM_MEM[3876] = 8'h9E;
ROM_MEM[3877] = 8'h19;
ROM_MEM[3878] = 8'hC7;
ROM_MEM[3879] = 8'h1C;
ROM_MEM[3880] = 8'h9D;
ROM_MEM[3881] = 8'h8B;
ROM_MEM[3882] = 8'h88;
ROM_MEM[3883] = 8'h85;
ROM_MEM[3884] = 8'hDD;
ROM_MEM[3885] = 8'h07;
ROM_MEM[3886] = 8'hFF;
ROM_MEM[3887] = 8'hFF;
ROM_MEM[3888] = 8'hFF;
ROM_MEM[3889] = 8'h04;
ROM_MEM[3890] = 8'h30;
ROM_MEM[3891] = 8'h3A;
ROM_MEM[3892] = 8'hBC;
ROM_MEM[3893] = 8'h2D;
ROM_MEM[3894] = 8'hD1;
ROM_MEM[3895] = 8'h17;
ROM_MEM[3896] = 8'hAB;
ROM_MEM[3897] = 8'h6E;
ROM_MEM[3898] = 8'h91;
ROM_MEM[3899] = 8'hB2;
ROM_MEM[3900] = 8'h07;
ROM_MEM[3901] = 8'h95;
ROM_MEM[3902] = 8'hA2;
ROM_MEM[3903] = 8'h1E;
ROM_MEM[3904] = 8'h49;
ROM_MEM[3905] = 8'h14;
ROM_MEM[3906] = 8'h60;
ROM_MEM[3907] = 8'h94;
ROM_MEM[3908] = 8'hAB;
ROM_MEM[3909] = 8'h02;
ROM_MEM[3910] = 8'hB2;
ROM_MEM[3911] = 8'h37;
ROM_MEM[3912] = 8'h33;
ROM_MEM[3913] = 8'h40;
ROM_MEM[3914] = 8'h4A;
ROM_MEM[3915] = 8'h65;
ROM_MEM[3916] = 8'h06;
ROM_MEM[3917] = 8'h60;
ROM_MEM[3918] = 8'h5B;
ROM_MEM[3919] = 8'h7C;
ROM_MEM[3920] = 8'hF5;
ROM_MEM[3921] = 8'h7E;
ROM_MEM[3922] = 8'h99;
ROM_MEM[3923] = 8'h68;
ROM_MEM[3924] = 8'h76;
ROM_MEM[3925] = 8'hE5;
ROM_MEM[3926] = 8'h35;
ROM_MEM[3927] = 8'hF8;
ROM_MEM[3928] = 8'h1E;
ROM_MEM[3929] = 8'h4E;
ROM_MEM[3930] = 8'h52;
ROM_MEM[3931] = 8'h93;
ROM_MEM[3932] = 8'hD7;
ROM_MEM[3933] = 8'hE0;
ROM_MEM[3934] = 8'h5B;
ROM_MEM[3935] = 8'h3A;
ROM_MEM[3936] = 8'h4B;
ROM_MEM[3937] = 8'h4C;
ROM_MEM[3938] = 8'h59;
ROM_MEM[3939] = 8'hA3;
ROM_MEM[3940] = 8'hAF;
ROM_MEM[3941] = 8'hE9;
ROM_MEM[3942] = 8'hAC;
ROM_MEM[3943] = 8'h31;
ROM_MEM[3944] = 8'h65;
ROM_MEM[3945] = 8'hCD;
ROM_MEM[3946] = 8'h61;
ROM_MEM[3947] = 8'h44;
ROM_MEM[3948] = 8'h90;
ROM_MEM[3949] = 8'hD6;
ROM_MEM[3950] = 8'h94;
ROM_MEM[3951] = 8'hB5;
ROM_MEM[3952] = 8'hC5;
ROM_MEM[3953] = 8'hE0;
ROM_MEM[3954] = 8'h4D;
ROM_MEM[3955] = 8'h5C;
ROM_MEM[3956] = 8'h95;
ROM_MEM[3957] = 8'hC7;
ROM_MEM[3958] = 8'h50;
ROM_MEM[3959] = 8'hC5;
ROM_MEM[3960] = 8'hBA;
ROM_MEM[3961] = 8'hA8;
ROM_MEM[3962] = 8'hC5;
ROM_MEM[3963] = 8'h4E;
ROM_MEM[3964] = 8'hC0;
ROM_MEM[3965] = 8'h02;
ROM_MEM[3966] = 8'h96;
ROM_MEM[3967] = 8'h09;
ROM_MEM[3968] = 8'h98;
ROM_MEM[3969] = 8'h24;
ROM_MEM[3970] = 8'h2B;
ROM_MEM[3971] = 8'h00;
ROM_MEM[3972] = 8'h55;
ROM_MEM[3973] = 8'h54;
ROM_MEM[3974] = 8'h29;
ROM_MEM[3975] = 8'h20;
ROM_MEM[3976] = 8'h8B;
ROM_MEM[3977] = 8'h52;
ROM_MEM[3978] = 8'h01;
ROM_MEM[3979] = 8'h24;
ROM_MEM[3980] = 8'h5E;
ROM_MEM[3981] = 8'h5A;
ROM_MEM[3982] = 8'h1A;
ROM_MEM[3983] = 8'hE7;
ROM_MEM[3984] = 8'h5B;
ROM_MEM[3985] = 8'hC5;
ROM_MEM[3986] = 8'hAA;
ROM_MEM[3987] = 8'h76;
ROM_MEM[3988] = 8'h9B;
ROM_MEM[3989] = 8'h43;
ROM_MEM[3990] = 8'hF4;
ROM_MEM[3991] = 8'h60;
ROM_MEM[3992] = 8'hAE;
ROM_MEM[3993] = 8'hC6;
ROM_MEM[3994] = 8'h6D;
ROM_MEM[3995] = 8'h09;
ROM_MEM[3996] = 8'hC9;
ROM_MEM[3997] = 8'h13;
ROM_MEM[3998] = 8'hB9;
ROM_MEM[3999] = 8'h1B;
ROM_MEM[4000] = 8'h97;
ROM_MEM[4001] = 8'hD5;
ROM_MEM[4002] = 8'h67;
ROM_MEM[4003] = 8'h37;
ROM_MEM[4004] = 8'h96;
ROM_MEM[4005] = 8'hAA;
ROM_MEM[4006] = 8'h5D;
ROM_MEM[4007] = 8'h56;
ROM_MEM[4008] = 8'hCD;
ROM_MEM[4009] = 8'h2B;
ROM_MEM[4010] = 8'hD2;
ROM_MEM[4011] = 8'h2C;
ROM_MEM[4012] = 8'h71;
ROM_MEM[4013] = 8'hD8;
ROM_MEM[4014] = 8'h3D;
ROM_MEM[4015] = 8'h8B;
ROM_MEM[4016] = 8'hCC;
ROM_MEM[4017] = 8'hF0;
ROM_MEM[4018] = 8'h24;
ROM_MEM[4019] = 8'h6D;
ROM_MEM[4020] = 8'h0A;
ROM_MEM[4021] = 8'h5E;
ROM_MEM[4022] = 8'hDC;
ROM_MEM[4023] = 8'h2A;
ROM_MEM[4024] = 8'h6B;
ROM_MEM[4025] = 8'h8F;
ROM_MEM[4026] = 8'h35;
ROM_MEM[4027] = 8'h38;
ROM_MEM[4028] = 8'h4E;
ROM_MEM[4029] = 8'hAF;
ROM_MEM[4030] = 8'hAC;
ROM_MEM[4031] = 8'hD5;
ROM_MEM[4032] = 8'h56;
ROM_MEM[4033] = 8'h1F;
ROM_MEM[4034] = 8'h39;
ROM_MEM[4035] = 8'hBC;
ROM_MEM[4036] = 8'hAA;
ROM_MEM[4037] = 8'h56;
ROM_MEM[4038] = 8'h59;
ROM_MEM[4039] = 8'h7D;
ROM_MEM[4040] = 8'hB0;
ROM_MEM[4041] = 8'h50;
ROM_MEM[4042] = 8'h8D;
ROM_MEM[4043] = 8'h46;
ROM_MEM[4044] = 8'h69;
ROM_MEM[4045] = 8'h37;
ROM_MEM[4046] = 8'h2E;
ROM_MEM[4047] = 8'hCC;
ROM_MEM[4048] = 8'hC5;
ROM_MEM[4049] = 8'h1A;
ROM_MEM[4050] = 8'h97;
ROM_MEM[4051] = 8'hD5;
ROM_MEM[4052] = 8'h67;
ROM_MEM[4053] = 8'h33;
ROM_MEM[4054] = 8'h95;
ROM_MEM[4055] = 8'h6C;
ROM_MEM[4056] = 8'hDC;
ROM_MEM[4057] = 8'h16;
ROM_MEM[4058] = 8'h9F;
ROM_MEM[4059] = 8'h25;
ROM_MEM[4060] = 8'h34;
ROM_MEM[4061] = 8'hAB;
ROM_MEM[4062] = 8'hF6;
ROM_MEM[4063] = 8'h58;
ROM_MEM[4064] = 8'h63;
ROM_MEM[4065] = 8'hA2;
ROM_MEM[4066] = 8'hB0;
ROM_MEM[4067] = 8'h9A;
ROM_MEM[4068] = 8'hC8;
ROM_MEM[4069] = 8'h63;
ROM_MEM[4070] = 8'h0B;
ROM_MEM[4071] = 8'h91;
ROM_MEM[4072] = 8'hAD;
ROM_MEM[4073] = 8'h62;
ROM_MEM[4074] = 8'hAC;
ROM_MEM[4075] = 8'h94;
ROM_MEM[4076] = 8'hC3;
ROM_MEM[4077] = 8'hEB;
ROM_MEM[4078] = 8'hD0;
ROM_MEM[4079] = 8'h88;
ROM_MEM[4080] = 8'hB2;
ROM_MEM[4081] = 8'h9D;
ROM_MEM[4082] = 8'hD6;
ROM_MEM[4083] = 8'h2C;
ROM_MEM[4084] = 8'h42;
ROM_MEM[4085] = 8'h3C;
ROM_MEM[4086] = 8'h2C;
ROM_MEM[4087] = 8'h4E;
ROM_MEM[4088] = 8'hF9;
ROM_MEM[4089] = 8'h82;
ROM_MEM[4090] = 8'h08;
ROM_MEM[4091] = 8'h8B;
ROM_MEM[4092] = 8'h2C;
ROM_MEM[4093] = 8'hDB;
ROM_MEM[4094] = 8'h0A;
ROM_MEM[4095] = 8'h80;
ROM_MEM[4096] = 8'h35;
ROM_MEM[4097] = 8'hB3;
ROM_MEM[4098] = 8'hFC;
ROM_MEM[4099] = 8'hDE;
ROM_MEM[4100] = 8'h4A;
ROM_MEM[4101] = 8'h74;
ROM_MEM[4102] = 8'hA5;
ROM_MEM[4103] = 8'h25;
ROM_MEM[4104] = 8'h03;
ROM_MEM[4105] = 8'hD0;
ROM_MEM[4106] = 8'h62;
ROM_MEM[4107] = 8'h5D;
ROM_MEM[4108] = 8'h5E;
ROM_MEM[4109] = 8'h13;
ROM_MEM[4110] = 8'h3C;
ROM_MEM[4111] = 8'h33;
ROM_MEM[4112] = 8'h2A;
ROM_MEM[4113] = 8'h52;
ROM_MEM[4114] = 8'hFA;
ROM_MEM[4115] = 8'hBC;
ROM_MEM[4116] = 8'h0D;
ROM_MEM[4117] = 8'h77;
ROM_MEM[4118] = 8'hCF;
ROM_MEM[4119] = 8'h84;
ROM_MEM[4120] = 8'hE1;
ROM_MEM[4121] = 8'h0F;
ROM_MEM[4122] = 8'hCA;
ROM_MEM[4123] = 8'hDD;
ROM_MEM[4124] = 8'hD5;
ROM_MEM[4125] = 8'h5B;
ROM_MEM[4126] = 8'h31;
ROM_MEM[4127] = 8'h40;
ROM_MEM[4128] = 8'h45;
ROM_MEM[4129] = 8'h13;
ROM_MEM[4130] = 8'h06;
ROM_MEM[4131] = 8'h98;
ROM_MEM[4132] = 8'hE2;
ROM_MEM[4133] = 8'h42;
ROM_MEM[4134] = 8'h00;
ROM_MEM[4135] = 8'hA3;
ROM_MEM[4136] = 8'hC3;
ROM_MEM[4137] = 8'hE0;
ROM_MEM[4138] = 8'h01;
ROM_MEM[4139] = 8'h00;
ROM_MEM[4140] = 8'h00;
ROM_MEM[4141] = 8'h00;
ROM_MEM[4142] = 8'h40;
ROM_MEM[4143] = 8'h80;
ROM_MEM[4144] = 8'h8C;
ROM_MEM[4145] = 8'h32;
ROM_MEM[4146] = 8'h08;
ROM_MEM[4147] = 8'h10;
ROM_MEM[4148] = 8'h6C;
ROM_MEM[4149] = 8'h06;
ROM_MEM[4150] = 8'h03;
ROM_MEM[4151] = 8'h7C;
ROM_MEM[4152] = 8'h2A;
ROM_MEM[4153] = 8'h69;
ROM_MEM[4154] = 8'h53;
ROM_MEM[4155] = 8'h08;
ROM_MEM[4156] = 8'hDD;
ROM_MEM[4157] = 8'h2C;
ROM_MEM[4158] = 8'h52;
ROM_MEM[4159] = 8'hA7;
ROM_MEM[4160] = 8'hAD;
ROM_MEM[4161] = 8'h7E;
ROM_MEM[4162] = 8'h56;
ROM_MEM[4163] = 8'hB0;
ROM_MEM[4164] = 8'h78;
ROM_MEM[4165] = 8'hA3;
ROM_MEM[4166] = 8'hB6;
ROM_MEM[4167] = 8'hFA;
ROM_MEM[4168] = 8'h95;
ROM_MEM[4169] = 8'hCE;
ROM_MEM[4170] = 8'h1A;
ROM_MEM[4171] = 8'hB3;
ROM_MEM[4172] = 8'hDA;
ROM_MEM[4173] = 8'hEA;
ROM_MEM[4174] = 8'h47;
ROM_MEM[4175] = 8'h24;
ROM_MEM[4176] = 8'h6B;
ROM_MEM[4177] = 8'hD6;
ROM_MEM[4178] = 8'h6E;
ROM_MEM[4179] = 8'h7B;
ROM_MEM[4180] = 8'h68;
ROM_MEM[4181] = 8'h19;
ROM_MEM[4182] = 8'hA8;
ROM_MEM[4183] = 8'hDE;
ROM_MEM[4184] = 8'hB8;
ROM_MEM[4185] = 8'h1D;
ROM_MEM[4186] = 8'h21;
ROM_MEM[4187] = 8'hF8;
ROM_MEM[4188] = 8'h30;
ROM_MEM[4189] = 8'h45;
ROM_MEM[4190] = 8'hEB;
ROM_MEM[4191] = 8'h74;
ROM_MEM[4192] = 8'hF8;
ROM_MEM[4193] = 8'h10;
ROM_MEM[4194] = 8'h69;
ROM_MEM[4195] = 8'h68;
ROM_MEM[4196] = 8'h8D;
ROM_MEM[4197] = 8'hD3;
ROM_MEM[4198] = 8'hE1;
ROM_MEM[4199] = 8'h4D;
ROM_MEM[4200] = 8'h87;
ROM_MEM[4201] = 8'hAB;
ROM_MEM[4202] = 8'h27;
ROM_MEM[4203] = 8'h16;
ROM_MEM[4204] = 8'h00;
ROM_MEM[4205] = 8'h6A;
ROM_MEM[4206] = 8'h29;
ROM_MEM[4207] = 8'hE5;
ROM_MEM[4208] = 8'hF3;
ROM_MEM[4209] = 8'hA1;
ROM_MEM[4210] = 8'h5C;
ROM_MEM[4211] = 8'hD5;
ROM_MEM[4212] = 8'h5B;
ROM_MEM[4213] = 8'h1B;
ROM_MEM[4214] = 8'h80;
ROM_MEM[4215] = 8'h26;
ROM_MEM[4216] = 8'hEB;
ROM_MEM[4217] = 8'hF6;
ROM_MEM[4218] = 8'hA7;
ROM_MEM[4219] = 8'h28;
ROM_MEM[4220] = 8'hA6;
ROM_MEM[4221] = 8'h9A;
ROM_MEM[4222] = 8'h21;
ROM_MEM[4223] = 8'h15;
ROM_MEM[4224] = 8'hC0;
ROM_MEM[4225] = 8'hB3;
ROM_MEM[4226] = 8'h95;
ROM_MEM[4227] = 8'h02;
ROM_MEM[4228] = 8'h68;
ROM_MEM[4229] = 8'hB5;
ROM_MEM[4230] = 8'h14;
ROM_MEM[4231] = 8'h80;
ROM_MEM[4232] = 8'h2F;
ROM_MEM[4233] = 8'h5A;
ROM_MEM[4234] = 8'h02;
ROM_MEM[4235] = 8'hF0;
ROM_MEM[4236] = 8'h21;
ROM_MEM[4237] = 8'hC2;
ROM_MEM[4238] = 8'h00;
ROM_MEM[4239] = 8'h95;
ROM_MEM[4240] = 8'hBA;
ROM_MEM[4241] = 8'h28;
ROM_MEM[4242] = 8'h60;
ROM_MEM[4243] = 8'h00;
ROM_MEM[4244] = 8'h33;
ROM_MEM[4245] = 8'h01;
ROM_MEM[4246] = 8'h1C;
ROM_MEM[4247] = 8'h24;
ROM_MEM[4248] = 8'h2E;
ROM_MEM[4249] = 8'h80;
ROM_MEM[4250] = 8'h8B;
ROM_MEM[4251] = 8'h25;
ROM_MEM[4252] = 8'h18;
ROM_MEM[4253] = 8'h90;
ROM_MEM[4254] = 8'hA1;
ROM_MEM[4255] = 8'h3B;
ROM_MEM[4256] = 8'h05;
ROM_MEM[4257] = 8'h30;
ROM_MEM[4258] = 8'hF0;
ROM_MEM[4259] = 8'h00;
ROM_MEM[4260] = 8'h9F;
ROM_MEM[4261] = 8'h0F;
ROM_MEM[4262] = 8'hE5;
ROM_MEM[4263] = 8'h0D;
ROM_MEM[4264] = 8'hAC;
ROM_MEM[4265] = 8'hC9;
ROM_MEM[4266] = 8'hCB;
ROM_MEM[4267] = 8'hC2;
ROM_MEM[4268] = 8'hE3;
ROM_MEM[4269] = 8'h1D;
ROM_MEM[4270] = 8'hA8;
ROM_MEM[4271] = 8'hC4;
ROM_MEM[4272] = 8'h68;
ROM_MEM[4273] = 8'hAB;
ROM_MEM[4274] = 8'h4C;
ROM_MEM[4275] = 8'h79;
ROM_MEM[4276] = 8'hB0;
ROM_MEM[4277] = 8'h96;
ROM_MEM[4278] = 8'hAB;
ROM_MEM[4279] = 8'h25;
ROM_MEM[4280] = 8'h2D;
ROM_MEM[4281] = 8'hD9;
ROM_MEM[4282] = 8'hC1;
ROM_MEM[4283] = 8'h47;
ROM_MEM[4284] = 8'hAF;
ROM_MEM[4285] = 8'hAC;
ROM_MEM[4286] = 8'hB0;
ROM_MEM[4287] = 8'h38;
ROM_MEM[4288] = 8'h47;
ROM_MEM[4289] = 8'hEC;
ROM_MEM[4290] = 8'hAD;
ROM_MEM[4291] = 8'h52;
ROM_MEM[4292] = 8'hCB;
ROM_MEM[4293] = 8'h92;
ROM_MEM[4294] = 8'h2C;
ROM_MEM[4295] = 8'hA9;
ROM_MEM[4296] = 8'hB5;
ROM_MEM[4297] = 8'h18;
ROM_MEM[4298] = 8'h6D;
ROM_MEM[4299] = 8'h8B;
ROM_MEM[4300] = 8'hEB;
ROM_MEM[4301] = 8'h80;
ROM_MEM[4302] = 8'h3A;
ROM_MEM[4303] = 8'h7C;
ROM_MEM[4304] = 8'h04;
ROM_MEM[4305] = 8'h10;
ROM_MEM[4306] = 8'h02;
ROM_MEM[4307] = 8'h38;
ROM_MEM[4308] = 8'h01;
ROM_MEM[4309] = 8'h00;
ROM_MEM[4310] = 8'h55;
ROM_MEM[4311] = 8'h25;
ROM_MEM[4312] = 8'h00;
ROM_MEM[4313] = 8'h40;
ROM_MEM[4314] = 8'h6A;
ROM_MEM[4315] = 8'h08;
ROM_MEM[4316] = 8'h00;
ROM_MEM[4317] = 8'h50;
ROM_MEM[4318] = 8'h8C;
ROM_MEM[4319] = 8'h00;
ROM_MEM[4320] = 8'h00;
ROM_MEM[4321] = 8'h89;
ROM_MEM[4322] = 8'h2B;
ROM_MEM[4323] = 8'hC0;
ROM_MEM[4324] = 8'h6A;
ROM_MEM[4325] = 8'h91;
ROM_MEM[4326] = 8'h05;
ROM_MEM[4327] = 8'hCC;
ROM_MEM[4328] = 8'hD6;
ROM_MEM[4329] = 8'hD3;
ROM_MEM[4330] = 8'hC0;
ROM_MEM[4331] = 8'h38;
ROM_MEM[4332] = 8'h63;
ROM_MEM[4333] = 8'h5D;
ROM_MEM[4334] = 8'hBA;
ROM_MEM[4335] = 8'h55;
ROM_MEM[4336] = 8'h01;
ROM_MEM[4337] = 8'hA3;
ROM_MEM[4338] = 8'hE5;
ROM_MEM[4339] = 8'hCB;
ROM_MEM[4340] = 8'h8C;
ROM_MEM[4341] = 8'h98;
ROM_MEM[4342] = 8'h85;
ROM_MEM[4343] = 8'h8C;
ROM_MEM[4344] = 8'hCC;
ROM_MEM[4345] = 8'h75;
ROM_MEM[4346] = 8'h5B;
ROM_MEM[4347] = 8'h93;
ROM_MEM[4348] = 8'h3A;
ROM_MEM[4349] = 8'hDE;
ROM_MEM[4350] = 8'hA3;
ROM_MEM[4351] = 8'h75;
ROM_MEM[4352] = 8'hE9;
ROM_MEM[4353] = 8'hB0;
ROM_MEM[4354] = 8'hEB;
ROM_MEM[4355] = 8'h24;
ROM_MEM[4356] = 8'h4F;
ROM_MEM[4357] = 8'h26;
ROM_MEM[4358] = 8'h24;
ROM_MEM[4359] = 8'hD3;
ROM_MEM[4360] = 8'hAE;
ROM_MEM[4361] = 8'h93;
ROM_MEM[4362] = 8'h3C;
ROM_MEM[4363] = 8'h19;
ROM_MEM[4364] = 8'h97;
ROM_MEM[4365] = 8'h2C;
ROM_MEM[4366] = 8'hAB;
ROM_MEM[4367] = 8'h4A;
ROM_MEM[4368] = 8'h8C;
ROM_MEM[4369] = 8'hCA;
ROM_MEM[4370] = 8'hC9;
ROM_MEM[4371] = 8'h3A;
ROM_MEM[4372] = 8'hED;
ROM_MEM[4373] = 8'h3A;
ROM_MEM[4374] = 8'hE0;
ROM_MEM[4375] = 8'h62;
ROM_MEM[4376] = 8'hC4;
ROM_MEM[4377] = 8'h00;
ROM_MEM[4378] = 8'hAC;
ROM_MEM[4379] = 8'hB7;
ROM_MEM[4380] = 8'hC7;
ROM_MEM[4381] = 8'h80;
ROM_MEM[4382] = 8'hF6;
ROM_MEM[4383] = 8'hFD;
ROM_MEM[4384] = 8'h0B;
ROM_MEM[4385] = 8'hB8;
ROM_MEM[4386] = 8'hFB;
ROM_MEM[4387] = 8'hD6;
ROM_MEM[4388] = 8'hFD;
ROM_MEM[4389] = 8'hDB;
ROM_MEM[4390] = 8'h6E;
ROM_MEM[4391] = 8'h60;
ROM_MEM[4392] = 8'h3A;
ROM_MEM[4393] = 8'hDE;
ROM_MEM[4394] = 8'h6E;
ROM_MEM[4395] = 8'h3B;
ROM_MEM[4396] = 8'hA7;
ROM_MEM[4397] = 8'h80;
ROM_MEM[4398] = 8'hD1;
ROM_MEM[4399] = 8'hC9;
ROM_MEM[4400] = 8'h65;
ROM_MEM[4401] = 8'h78;
ROM_MEM[4402] = 8'hA4;
ROM_MEM[4403] = 8'h82;
ROM_MEM[4404] = 8'h27;
ROM_MEM[4405] = 8'hC5;
ROM_MEM[4406] = 8'hFA;
ROM_MEM[4407] = 8'h69;
ROM_MEM[4408] = 8'h49;
ROM_MEM[4409] = 8'hCA;
ROM_MEM[4410] = 8'h1E;
ROM_MEM[4411] = 8'hD0;
ROM_MEM[4412] = 8'h84;
ROM_MEM[4413] = 8'h74;
ROM_MEM[4414] = 8'hC4;
ROM_MEM[4415] = 8'h09;
ROM_MEM[4416] = 8'hB9;
ROM_MEM[4417] = 8'h23;
ROM_MEM[4418] = 8'hEB;
ROM_MEM[4419] = 8'h52;
ROM_MEM[4420] = 8'h61;
ROM_MEM[4421] = 8'h27;
ROM_MEM[4422] = 8'hE4;
ROM_MEM[4423] = 8'h9E;
ROM_MEM[4424] = 8'h8C;
ROM_MEM[4425] = 8'h4B;
ROM_MEM[4426] = 8'h86;
ROM_MEM[4427] = 8'h5D;
ROM_MEM[4428] = 8'h23;
ROM_MEM[4429] = 8'h19;
ROM_MEM[4430] = 8'h31;
ROM_MEM[4431] = 8'h6E;
ROM_MEM[4432] = 8'h19;
ROM_MEM[4433] = 8'h76;
ROM_MEM[4434] = 8'h03;
ROM_MEM[4435] = 8'hB0;
ROM_MEM[4436] = 8'h19;
ROM_MEM[4437] = 8'h62;
ROM_MEM[4438] = 8'h08;
ROM_MEM[4439] = 8'hF7;
ROM_MEM[4440] = 8'hBB;
ROM_MEM[4441] = 8'hEB;
ROM_MEM[4442] = 8'h7F;
ROM_MEM[4443] = 8'hDB;
ROM_MEM[4444] = 8'h0E;
ROM_MEM[4445] = 8'hE8;
ROM_MEM[4446] = 8'h3F;
ROM_MEM[4447] = 8'h2E;
ROM_MEM[4448] = 8'h80;
ROM_MEM[4449] = 8'hF1;
ROM_MEM[4450] = 8'hA7;
ROM_MEM[4451] = 8'hDB;
ROM_MEM[4452] = 8'h6E;
ROM_MEM[4453] = 8'h1C;
ROM_MEM[4454] = 8'h03;
ROM_MEM[4455] = 8'hFA;
ROM_MEM[4456] = 8'h5F;
ROM_MEM[4457] = 8'hA5;
ROM_MEM[4458] = 8'h32;
ROM_MEM[4459] = 8'h6B;
ROM_MEM[4460] = 8'h42;
ROM_MEM[4461] = 8'hE7;
ROM_MEM[4462] = 8'h7F;
ROM_MEM[4463] = 8'h95;
ROM_MEM[4464] = 8'h73;
ROM_MEM[4465] = 8'hAE;
ROM_MEM[4466] = 8'hCD;
ROM_MEM[4467] = 8'h5D;
ROM_MEM[4468] = 8'hEA;
ROM_MEM[4469] = 8'hFC;
ROM_MEM[4470] = 8'hCF;
ROM_MEM[4471] = 8'h32;
ROM_MEM[4472] = 8'hA9;
ROM_MEM[4473] = 8'h35;
ROM_MEM[4474] = 8'hA1;
ROM_MEM[4475] = 8'hF3;
ROM_MEM[4476] = 8'hBF;
ROM_MEM[4477] = 8'hCA;
ROM_MEM[4478] = 8'h39;
ROM_MEM[4479] = 8'hD7;
ROM_MEM[4480] = 8'hA6;
ROM_MEM[4481] = 8'hCE;
ROM_MEM[4482] = 8'hFF;
ROM_MEM[4483] = 8'h4A;
ROM_MEM[4484] = 8'hE3;
ROM_MEM[4485] = 8'h5A;
ROM_MEM[4486] = 8'h1B;
ROM_MEM[4487] = 8'h3A;
ROM_MEM[4488] = 8'hFF;
ROM_MEM[4489] = 8'hAB;
ROM_MEM[4490] = 8'h8C;
ROM_MEM[4491] = 8'h6B;
ROM_MEM[4492] = 8'h6D;
ROM_MEM[4493] = 8'hEA;
ROM_MEM[4494] = 8'hFC;
ROM_MEM[4495] = 8'hEF;
ROM_MEM[4496] = 8'h74;
ROM_MEM[4497] = 8'hCE;
ROM_MEM[4498] = 8'hB5;
ROM_MEM[4499] = 8'hA9;
ROM_MEM[4500] = 8'hF3;
ROM_MEM[4501] = 8'hBF;
ROM_MEM[4502] = 8'hD2;
ROM_MEM[4503] = 8'hA5;
ROM_MEM[4504] = 8'hD6;
ROM_MEM[4505] = 8'hA6;
ROM_MEM[4506] = 8'hCE;
ROM_MEM[4507] = 8'hFF;
ROM_MEM[4508] = 8'h4A;
ROM_MEM[4509] = 8'h93;
ROM_MEM[4510] = 8'h5A;
ROM_MEM[4511] = 8'hFB;
ROM_MEM[4512] = 8'h00;
ROM_MEM[4513] = 8'hEB;
ROM_MEM[4514] = 8'h24;
ROM_MEM[4515] = 8'h4F;
ROM_MEM[4516] = 8'h0C;
ROM_MEM[4517] = 8'h30;
ROM_MEM[4518] = 8'h7D;
ROM_MEM[4519] = 8'h4A;
ROM_MEM[4520] = 8'h01;
ROM_MEM[4521] = 8'hB6;
ROM_MEM[4522] = 8'h54;
ROM_MEM[4523] = 8'h19;
ROM_MEM[4524] = 8'hC0;
ROM_MEM[4525] = 8'hB5;
ROM_MEM[4526] = 8'hAC;
ROM_MEM[4527] = 8'h84;
ROM_MEM[4528] = 8'h47;
ROM_MEM[4529] = 8'h63;
ROM_MEM[4530] = 8'h1D;
ROM_MEM[4531] = 8'hC9;
ROM_MEM[4532] = 8'h72;
ROM_MEM[4533] = 8'h02;
ROM_MEM[4534] = 8'h11;
ROM_MEM[4535] = 8'h6C;
ROM_MEM[4536] = 8'h64;
ROM_MEM[4537] = 8'h9A;
ROM_MEM[4538] = 8'h28;
ROM_MEM[4539] = 8'h4D;
ROM_MEM[4540] = 8'h78;
ROM_MEM[4541] = 8'h32;
ROM_MEM[4542] = 8'h92;
ROM_MEM[4543] = 8'hA5;
ROM_MEM[4544] = 8'hEA;
ROM_MEM[4545] = 8'h3A;
ROM_MEM[4546] = 8'hE1;
ROM_MEM[4547] = 8'hD9;
ROM_MEM[4548] = 8'hA8;
ROM_MEM[4549] = 8'h8C;
ROM_MEM[4550] = 8'hB9;
ROM_MEM[4551] = 8'h9D;
ROM_MEM[4552] = 8'h82;
ROM_MEM[4553] = 8'h07;
ROM_MEM[4554] = 8'hE3;
ROM_MEM[4555] = 8'h55;
ROM_MEM[4556] = 8'h6C;
ROM_MEM[4557] = 8'h4E;
ROM_MEM[4558] = 8'h1B;
ROM_MEM[4559] = 8'h1E;
ROM_MEM[4560] = 8'h94;
ROM_MEM[4561] = 8'h67;
ROM_MEM[4562] = 8'h85;
ROM_MEM[4563] = 8'h5B;
ROM_MEM[4564] = 8'h6D;
ROM_MEM[4565] = 8'h78;
ROM_MEM[4566] = 8'hD2;
ROM_MEM[4567] = 8'h5A;
ROM_MEM[4568] = 8'hA9;
ROM_MEM[4569] = 8'h6E;
ROM_MEM[4570] = 8'h37;
ROM_MEM[4571] = 8'h01;
ROM_MEM[4572] = 8'h3A;
ROM_MEM[4573] = 8'hFA;
ROM_MEM[4574] = 8'h34;
ROM_MEM[4575] = 8'h3C;
ROM_MEM[4576] = 8'hE8;
ROM_MEM[4577] = 8'h88;
ROM_MEM[4578] = 8'h2A;
ROM_MEM[4579] = 8'h93;
ROM_MEM[4580] = 8'h9B;
ROM_MEM[4581] = 8'h00;
ROM_MEM[4582] = 8'h53;
ROM_MEM[4583] = 8'h23;
ROM_MEM[4584] = 8'h13;
ROM_MEM[4585] = 8'h60;
ROM_MEM[4586] = 8'h72;
ROM_MEM[4587] = 8'h54;
ROM_MEM[4588] = 8'h23;
ROM_MEM[4589] = 8'hA2;
ROM_MEM[4590] = 8'hD6;
ROM_MEM[4591] = 8'h4A;
ROM_MEM[4592] = 8'h77;
ROM_MEM[4593] = 8'h29;
ROM_MEM[4594] = 8'h01;
ROM_MEM[4595] = 8'h10;
ROM_MEM[4596] = 8'h25;
ROM_MEM[4597] = 8'h2A;
ROM_MEM[4598] = 8'h00;
ROM_MEM[4599] = 8'hAE;
ROM_MEM[4600] = 8'h7B;
ROM_MEM[4601] = 8'h37;
ROM_MEM[4602] = 8'h32;
ROM_MEM[4603] = 8'h19;
ROM_MEM[4604] = 8'hF7;
ROM_MEM[4605] = 8'h4A;
ROM_MEM[4606] = 8'h13;
ROM_MEM[4607] = 8'h9B;
ROM_MEM[4608] = 8'h00;
ROM_MEM[4609] = 8'h3B;
ROM_MEM[4610] = 8'h32;
ROM_MEM[4611] = 8'h02;
ROM_MEM[4612] = 8'hE0;
ROM_MEM[4613] = 8'hA2;
ROM_MEM[4614] = 8'h67;
ROM_MEM[4615] = 8'h00;
ROM_MEM[4616] = 8'h6C;
ROM_MEM[4617] = 8'hF0;
ROM_MEM[4618] = 8'h2C;
ROM_MEM[4619] = 8'h64;
ROM_MEM[4620] = 8'h36;
ROM_MEM[4621] = 8'hAA;
ROM_MEM[4622] = 8'h15;
ROM_MEM[4623] = 8'h61;
ROM_MEM[4624] = 8'hB9;
ROM_MEM[4625] = 8'h91;
ROM_MEM[4626] = 8'hC9;
ROM_MEM[4627] = 8'h6A;
ROM_MEM[4628] = 8'h74;
ROM_MEM[4629] = 8'h98;
ROM_MEM[4630] = 8'hD4;
ROM_MEM[4631] = 8'h00;
ROM_MEM[4632] = 8'hB8;
ROM_MEM[4633] = 8'hE8;
ROM_MEM[4634] = 8'h9D;
ROM_MEM[4635] = 8'h00;
ROM_MEM[4636] = 8'h93;
ROM_MEM[4637] = 8'hA3;
ROM_MEM[4638] = 8'h1A;
ROM_MEM[4639] = 8'h99;
ROM_MEM[4640] = 8'h94;
ROM_MEM[4641] = 8'h47;
ROM_MEM[4642] = 8'h84;
ROM_MEM[4643] = 8'hDB;
ROM_MEM[4644] = 8'h09;
ROM_MEM[4645] = 8'h80;
ROM_MEM[4646] = 8'h29;
ROM_MEM[4647] = 8'h11;
ROM_MEM[4648] = 8'h85;
ROM_MEM[4649] = 8'h8C;
ROM_MEM[4650] = 8'h3A;
ROM_MEM[4651] = 8'hBC;
ROM_MEM[4652] = 8'hDC;
ROM_MEM[4653] = 8'hE4;
ROM_MEM[4654] = 8'h14;
ROM_MEM[4655] = 8'h32;
ROM_MEM[4656] = 8'h19;
ROM_MEM[4657] = 8'h8F;
ROM_MEM[4658] = 8'h0A;
ROM_MEM[4659] = 8'h95;
ROM_MEM[4660] = 8'hD2;
ROM_MEM[4661] = 8'hC8;
ROM_MEM[4662] = 8'h64;
ROM_MEM[4663] = 8'hC3;
ROM_MEM[4664] = 8'hA7;
ROM_MEM[4665] = 8'h54;
ROM_MEM[4666] = 8'h6E;
ROM_MEM[4667] = 8'h21;
ROM_MEM[4668] = 8'hA3;
ROM_MEM[4669] = 8'h4A;
ROM_MEM[4670] = 8'h8F;
ROM_MEM[4671] = 8'h54;
ROM_MEM[4672] = 8'h3B;
ROM_MEM[4673] = 8'h01;
ROM_MEM[4674] = 8'h30;
ROM_MEM[4675] = 8'h35;
ROM_MEM[4676] = 8'h2A;
ROM_MEM[4677] = 8'h00;
ROM_MEM[4678] = 8'h2E;
ROM_MEM[4679] = 8'h45;
ROM_MEM[4680] = 8'h06;
ROM_MEM[4681] = 8'hC0;
ROM_MEM[4682] = 8'hC6;
ROM_MEM[4683] = 8'hF2;
ROM_MEM[4684] = 8'h42;
ROM_MEM[4685] = 8'h27;
ROM_MEM[4686] = 8'h13;
ROM_MEM[4687] = 8'h99;
ROM_MEM[4688] = 8'h13;
ROM_MEM[4689] = 8'hF4;
ROM_MEM[4690] = 8'h1C;
ROM_MEM[4691] = 8'hE0;
ROM_MEM[4692] = 8'h63;
ROM_MEM[4693] = 8'h64;
ROM_MEM[4694] = 8'hA1;
ROM_MEM[4695] = 8'hB2;
ROM_MEM[4696] = 8'hF6;
ROM_MEM[4697] = 8'h88;
ROM_MEM[4698] = 8'h32;
ROM_MEM[4699] = 8'h39;
ROM_MEM[4700] = 8'h01;
ROM_MEM[4701] = 8'h30;
ROM_MEM[4702] = 8'h25;
ROM_MEM[4703] = 8'h32;
ROM_MEM[4704] = 8'h00;
ROM_MEM[4705] = 8'hA6;
ROM_MEM[4706] = 8'h44;
ROM_MEM[4707] = 8'h39;
ROM_MEM[4708] = 8'hC0;
ROM_MEM[4709] = 8'h96;
ROM_MEM[4710] = 8'hCA;
ROM_MEM[4711] = 8'h00;
ROM_MEM[4712] = 8'hB8;
ROM_MEM[4713] = 8'h52;
ROM_MEM[4714] = 8'hE5;
ROM_MEM[4715] = 8'h00;
ROM_MEM[4716] = 8'h9F;
ROM_MEM[4717] = 8'hAB;
ROM_MEM[4718] = 8'h0A;
ROM_MEM[4719] = 8'h15;
ROM_MEM[4720] = 8'h7C;
ROM_MEM[4721] = 8'hD6;
ROM_MEM[4722] = 8'h4C;
ROM_MEM[4723] = 8'hDA;
ROM_MEM[4724] = 8'h71;
ROM_MEM[4725] = 8'h80;
ROM_MEM[4726] = 8'h99;
ROM_MEM[4727] = 8'hD1;
ROM_MEM[4728] = 8'h0E;
ROM_MEM[4729] = 8'h30;
ROM_MEM[4730] = 8'hBB;
ROM_MEM[4731] = 8'hCA;
ROM_MEM[4732] = 8'h01;
ROM_MEM[4733] = 8'hFA;
ROM_MEM[4734] = 8'h46;
ROM_MEM[4735] = 8'h1B;
ROM_MEM[4736] = 8'h40;
ROM_MEM[4737] = 8'h5E;
ROM_MEM[4738] = 8'h4F;
ROM_MEM[4739] = 8'h05;
ROM_MEM[4740] = 8'hE8;
ROM_MEM[4741] = 8'h17;
ROM_MEM[4742] = 8'h29;
ROM_MEM[4743] = 8'h00;
ROM_MEM[4744] = 8'hB5;
ROM_MEM[4745] = 8'h23;
ROM_MEM[4746] = 8'h04;
ROM_MEM[4747] = 8'h20;
ROM_MEM[4748] = 8'h67;
ROM_MEM[4749] = 8'hB8;
ROM_MEM[4750] = 8'h00;
ROM_MEM[4751] = 8'hE4;
ROM_MEM[4752] = 8'hF0;
ROM_MEM[4753] = 8'h10;
ROM_MEM[4754] = 8'h80;
ROM_MEM[4755] = 8'hAE;
ROM_MEM[4756] = 8'h1E;
ROM_MEM[4757] = 8'h02;
ROM_MEM[4758] = 8'hD0;
ROM_MEM[4759] = 8'h35;
ROM_MEM[4760] = 8'h9D;
ROM_MEM[4761] = 8'h01;
ROM_MEM[4762] = 8'hA6;
ROM_MEM[4763] = 8'h95;
ROM_MEM[4764] = 8'h33;
ROM_MEM[4765] = 8'hC0;
ROM_MEM[4766] = 8'hD4;
ROM_MEM[4767] = 8'h74;
ROM_MEM[4768] = 8'h02;
ROM_MEM[4769] = 8'h98;
ROM_MEM[4770] = 8'h98;
ROM_MEM[4771] = 8'hCE;
ROM_MEM[4772] = 8'h00;
ROM_MEM[4773] = 8'h16;
ROM_MEM[4774] = 8'hCB;
ROM_MEM[4775] = 8'h19;
ROM_MEM[4776] = 8'h20;
ROM_MEM[4777] = 8'h53;
ROM_MEM[4778] = 8'h3A;
ROM_MEM[4779] = 8'h01;
ROM_MEM[4780] = 8'h4C;
ROM_MEM[4781] = 8'hC8;
ROM_MEM[4782] = 8'h20;
ROM_MEM[4783] = 8'h00;
ROM_MEM[4784] = 8'h4B;
ROM_MEM[4785] = 8'hE5;
ROM_MEM[4786] = 8'h04;
ROM_MEM[4787] = 8'h10;
ROM_MEM[4788] = 8'hA1;
ROM_MEM[4789] = 8'h82;
ROM_MEM[4790] = 8'h00;
ROM_MEM[4791] = 8'h2A;
ROM_MEM[4792] = 8'h96;
ROM_MEM[4793] = 8'h13;
ROM_MEM[4794] = 8'h20;
ROM_MEM[4795] = 8'hB8;
ROM_MEM[4796] = 8'h08;
ROM_MEM[4797] = 8'h04;
ROM_MEM[4798] = 8'h88;
ROM_MEM[4799] = 8'hD8;
ROM_MEM[4800] = 8'h41;
ROM_MEM[4801] = 8'h00;
ROM_MEM[4802] = 8'h65;
ROM_MEM[4803] = 8'h2B;
ROM_MEM[4804] = 8'h1E;
ROM_MEM[4805] = 8'h00;
ROM_MEM[4806] = 8'h87;
ROM_MEM[4807] = 8'h59;
ROM_MEM[4808] = 8'hC5;
ROM_MEM[4809] = 8'h48;
ROM_MEM[4810] = 8'h5B;
ROM_MEM[4811] = 8'h53;
ROM_MEM[4812] = 8'hB3;
ROM_MEM[4813] = 8'h6C;
ROM_MEM[4814] = 8'h2F;
ROM_MEM[4815] = 8'h2D;
ROM_MEM[4816] = 8'h4F;
ROM_MEM[4817] = 8'h2D;
ROM_MEM[4818] = 8'h1B;
ROM_MEM[4819] = 8'h97;
ROM_MEM[4820] = 8'hBD;
ROM_MEM[4821] = 8'hD4;
ROM_MEM[4822] = 8'h5A;
ROM_MEM[4823] = 8'h25;
ROM_MEM[4824] = 8'h78;
ROM_MEM[4825] = 8'hD5;
ROM_MEM[4826] = 8'h4E;
ROM_MEM[4827] = 8'h52;
ROM_MEM[4828] = 8'h7C;
ROM_MEM[4829] = 8'h34;
ROM_MEM[4830] = 8'hD3;
ROM_MEM[4831] = 8'h8C;
ROM_MEM[4832] = 8'hC8;
ROM_MEM[4833] = 8'h49;
ROM_MEM[4834] = 8'hF6;
ROM_MEM[4835] = 8'hC1;
ROM_MEM[4836] = 8'hCC;
ROM_MEM[4837] = 8'hCA;
ROM_MEM[4838] = 8'h2D;
ROM_MEM[4839] = 8'h36;
ROM_MEM[4840] = 8'h35;
ROM_MEM[4841] = 8'h07;
ROM_MEM[4842] = 8'hAC;
ROM_MEM[4843] = 8'h68;
ROM_MEM[4844] = 8'h91;
ROM_MEM[4845] = 8'h35;
ROM_MEM[4846] = 8'hE4;
ROM_MEM[4847] = 8'hE2;
ROM_MEM[4848] = 8'hB0;
ROM_MEM[4849] = 8'h32;
ROM_MEM[4850] = 8'h55;
ROM_MEM[4851] = 8'hD1;
ROM_MEM[4852] = 8'h10;
ROM_MEM[4853] = 8'hB3;
ROM_MEM[4854] = 8'hE5;
ROM_MEM[4855] = 8'hF6;
ROM_MEM[4856] = 8'h24;
ROM_MEM[4857] = 8'hC5;
ROM_MEM[4858] = 8'h83;
ROM_MEM[4859] = 8'h8F;
ROM_MEM[4860] = 8'h5E;
ROM_MEM[4861] = 8'hD6;
ROM_MEM[4862] = 8'h4D;
ROM_MEM[4863] = 8'h14;
ROM_MEM[4864] = 8'h1F;
ROM_MEM[4865] = 8'h36;
ROM_MEM[4866] = 8'h39;
ROM_MEM[4867] = 8'h9D;
ROM_MEM[4868] = 8'hDA;
ROM_MEM[4869] = 8'h60;
ROM_MEM[4870] = 8'h74;
ROM_MEM[4871] = 8'hE8;
ROM_MEM[4872] = 8'h64;
ROM_MEM[4873] = 8'h65;
ROM_MEM[4874] = 8'hB6;
ROM_MEM[4875] = 8'h43;
ROM_MEM[4876] = 8'h6B;
ROM_MEM[4877] = 8'hE3;
ROM_MEM[4878] = 8'hB3;
ROM_MEM[4879] = 8'hA5;
ROM_MEM[4880] = 8'hEA;
ROM_MEM[4881] = 8'h6B;
ROM_MEM[4882] = 8'hC5;
ROM_MEM[4883] = 8'hCE;
ROM_MEM[4884] = 8'h48;
ROM_MEM[4885] = 8'h5A;
ROM_MEM[4886] = 8'h22;
ROM_MEM[4887] = 8'h32;
ROM_MEM[4888] = 8'h24;
ROM_MEM[4889] = 8'hB9;
ROM_MEM[4890] = 8'h20;
ROM_MEM[4891] = 8'h69;
ROM_MEM[4892] = 8'hCD;
ROM_MEM[4893] = 8'h0A;
ROM_MEM[4894] = 8'hB3;
ROM_MEM[4895] = 8'hC4;
ROM_MEM[4896] = 8'h00;
ROM_MEM[4897] = 8'h17;
ROM_MEM[4898] = 8'hA2;
ROM_MEM[4899] = 8'h8A;
ROM_MEM[4900] = 8'h90;
ROM_MEM[4901] = 8'h2A;
ROM_MEM[4902] = 8'h85;
ROM_MEM[4903] = 8'h79;
ROM_MEM[4904] = 8'h59;
ROM_MEM[4905] = 8'h1E;
ROM_MEM[4906] = 8'h42;
ROM_MEM[4907] = 8'h74;
ROM_MEM[4908] = 8'hDA;
ROM_MEM[4909] = 8'h76;
ROM_MEM[4910] = 8'hE1;
ROM_MEM[4911] = 8'h38;
ROM_MEM[4912] = 8'hE8;
ROM_MEM[4913] = 8'h41;
ROM_MEM[4914] = 8'h4A;
ROM_MEM[4915] = 8'hA6;
ROM_MEM[4916] = 8'h87;
ROM_MEM[4917] = 8'h2C;
ROM_MEM[4918] = 8'hE7;
ROM_MEM[4919] = 8'h66;
ROM_MEM[4920] = 8'h65;
ROM_MEM[4921] = 8'h66;
ROM_MEM[4922] = 8'h91;
ROM_MEM[4923] = 8'h96;
ROM_MEM[4924] = 8'h8C;
ROM_MEM[4925] = 8'h96;
ROM_MEM[4926] = 8'hA4;
ROM_MEM[4927] = 8'h47;
ROM_MEM[4928] = 8'hA5;
ROM_MEM[4929] = 8'hD9;
ROM_MEM[4930] = 8'h0A;
ROM_MEM[4931] = 8'hBC;
ROM_MEM[4932] = 8'h73;
ROM_MEM[4933] = 8'hD9;
ROM_MEM[4934] = 8'h66;
ROM_MEM[4935] = 8'h21;
ROM_MEM[4936] = 8'h69;
ROM_MEM[4937] = 8'hB1;
ROM_MEM[4938] = 8'h29;
ROM_MEM[4939] = 8'h59;
ROM_MEM[4940] = 8'h68;
ROM_MEM[4941] = 8'hAD;
ROM_MEM[4942] = 8'hED;
ROM_MEM[4943] = 8'hC5;
ROM_MEM[4944] = 8'hA6;
ROM_MEM[4945] = 8'h16;
ROM_MEM[4946] = 8'h45;
ROM_MEM[4947] = 8'h9D;
ROM_MEM[4948] = 8'h72;
ROM_MEM[4949] = 8'h17;
ROM_MEM[4950] = 8'h9F;
ROM_MEM[4951] = 8'h9E;
ROM_MEM[4952] = 8'h59;
ROM_MEM[4953] = 8'h47;
ROM_MEM[4954] = 8'hC8;
ROM_MEM[4955] = 8'h59;
ROM_MEM[4956] = 8'h7C;
ROM_MEM[4957] = 8'h7A;
ROM_MEM[4958] = 8'hE6;
ROM_MEM[4959] = 8'h59;
ROM_MEM[4960] = 8'hED;
ROM_MEM[4961] = 8'h64;
ROM_MEM[4962] = 8'h09;
ROM_MEM[4963] = 8'h31;
ROM_MEM[4964] = 8'h47;
ROM_MEM[4965] = 8'h79;
ROM_MEM[4966] = 8'h37;
ROM_MEM[4967] = 8'h93;
ROM_MEM[4968] = 8'h60;
ROM_MEM[4969] = 8'h04;
ROM_MEM[4970] = 8'h6B;
ROM_MEM[4971] = 8'hCE;
ROM_MEM[4972] = 8'h19;
ROM_MEM[4973] = 8'hB2;
ROM_MEM[4974] = 8'h9D;
ROM_MEM[4975] = 8'h9B;
ROM_MEM[4976] = 8'hA2;
ROM_MEM[4977] = 8'h8B;
ROM_MEM[4978] = 8'hA8;
ROM_MEM[4979] = 8'hDA;
ROM_MEM[4980] = 8'h26;
ROM_MEM[4981] = 8'h40;
ROM_MEM[4982] = 8'h8C;
ROM_MEM[4983] = 8'hA6;
ROM_MEM[4984] = 8'h04;
ROM_MEM[4985] = 8'h08;
ROM_MEM[4986] = 8'hDA;
ROM_MEM[4987] = 8'hBD;
ROM_MEM[4988] = 8'hB0;
ROM_MEM[4989] = 8'h31;
ROM_MEM[4990] = 8'h4A;
ROM_MEM[4991] = 8'h57;
ROM_MEM[4992] = 8'hB6;
ROM_MEM[4993] = 8'h98;
ROM_MEM[4994] = 8'hC5;
ROM_MEM[4995] = 8'hA6;
ROM_MEM[4996] = 8'h20;
ROM_MEM[4997] = 8'h15;
ROM_MEM[4998] = 8'hD3;
ROM_MEM[4999] = 8'h4C;
ROM_MEM[5000] = 8'h0F;
ROM_MEM[5001] = 8'h97;
ROM_MEM[5002] = 8'h82;
ROM_MEM[5003] = 8'hD7;
ROM_MEM[5004] = 8'h78;
ROM_MEM[5005] = 8'hD2;
ROM_MEM[5006] = 8'h39;
ROM_MEM[5007] = 8'h7C;
ROM_MEM[5008] = 8'h89;
ROM_MEM[5009] = 8'h32;
ROM_MEM[5010] = 8'hB5;
ROM_MEM[5011] = 8'hE5;
ROM_MEM[5012] = 8'hE8;
ROM_MEM[5013] = 8'h08;
ROM_MEM[5014] = 8'h25;
ROM_MEM[5015] = 8'h6A;
ROM_MEM[5016] = 8'hC7;
ROM_MEM[5017] = 8'hA6;
ROM_MEM[5018] = 8'hDB;
ROM_MEM[5019] = 8'h23;
ROM_MEM[5020] = 8'h96;
ROM_MEM[5021] = 8'hA4;
ROM_MEM[5022] = 8'h95;
ROM_MEM[5023] = 8'h95;
ROM_MEM[5024] = 8'h6A;
ROM_MEM[5025] = 8'h8E;
ROM_MEM[5026] = 8'h9C;
ROM_MEM[5027] = 8'h53;
ROM_MEM[5028] = 8'h4C;
ROM_MEM[5029] = 8'h76;
ROM_MEM[5030] = 8'h32;
ROM_MEM[5031] = 8'h3D;
ROM_MEM[5032] = 8'h52;
ROM_MEM[5033] = 8'hF6;
ROM_MEM[5034] = 8'h36;
ROM_MEM[5035] = 8'hD1;
ROM_MEM[5036] = 8'hAE;
ROM_MEM[5037] = 8'h66;
ROM_MEM[5038] = 8'hB0;
ROM_MEM[5039] = 8'h29;
ROM_MEM[5040] = 8'h6A;
ROM_MEM[5041] = 8'hE9;
ROM_MEM[5042] = 8'hBA;
ROM_MEM[5043] = 8'hEB;
ROM_MEM[5044] = 8'hC5;
ROM_MEM[5045] = 8'hA6;
ROM_MEM[5046] = 8'h6E;
ROM_MEM[5047] = 8'hE9;
ROM_MEM[5048] = 8'hD5;
ROM_MEM[5049] = 8'hB2;
ROM_MEM[5050] = 8'h17;
ROM_MEM[5051] = 8'h13;
ROM_MEM[5052] = 8'h77;
ROM_MEM[5053] = 8'hBA;
ROM_MEM[5054] = 8'h45;
ROM_MEM[5055] = 8'h4B;
ROM_MEM[5056] = 8'h19;
ROM_MEM[5057] = 8'h4C;
ROM_MEM[5058] = 8'h78;
ROM_MEM[5059] = 8'h9E;
ROM_MEM[5060] = 8'h9A;
ROM_MEM[5061] = 8'h25;
ROM_MEM[5062] = 8'h65;
ROM_MEM[5063] = 8'hD0;
ROM_MEM[5064] = 8'hF1;
ROM_MEM[5065] = 8'h69;
ROM_MEM[5066] = 8'h44;
ROM_MEM[5067] = 8'h64;
ROM_MEM[5068] = 8'h94;
ROM_MEM[5069] = 8'h41;
ROM_MEM[5070] = 8'hC7;
ROM_MEM[5071] = 8'h2E;
ROM_MEM[5072] = 8'h2D;
ROM_MEM[5073] = 8'h3E;
ROM_MEM[5074] = 8'h4E;
ROM_MEM[5075] = 8'h1B;
ROM_MEM[5076] = 8'h1B;
ROM_MEM[5077] = 8'h0B;
ROM_MEM[5078] = 8'h4E;
ROM_MEM[5079] = 8'hC5;
ROM_MEM[5080] = 8'h24;
ROM_MEM[5081] = 8'h0E;
ROM_MEM[5082] = 8'h52;
ROM_MEM[5083] = 8'h08;
ROM_MEM[5084] = 8'hA6;
ROM_MEM[5085] = 8'h1E;
ROM_MEM[5086] = 8'h6A;
ROM_MEM[5087] = 8'h9B;
ROM_MEM[5088] = 8'h01;
ROM_MEM[5089] = 8'h71;
ROM_MEM[5090] = 8'h8A;
ROM_MEM[5091] = 8'h29;
ROM_MEM[5092] = 8'h20;
ROM_MEM[5093] = 8'hC5;
ROM_MEM[5094] = 8'h88;
ROM_MEM[5095] = 8'h42;
ROM_MEM[5096] = 8'h7B;
ROM_MEM[5097] = 8'hAB;
ROM_MEM[5098] = 8'hD9;
ROM_MEM[5099] = 8'hAE;
ROM_MEM[5100] = 8'h4A;
ROM_MEM[5101] = 8'h1B;
ROM_MEM[5102] = 8'hEB;
ROM_MEM[5103] = 8'hAD;
ROM_MEM[5104] = 8'hB6;
ROM_MEM[5105] = 8'h65;
ROM_MEM[5106] = 8'h52;
ROM_MEM[5107] = 8'h69;
ROM_MEM[5108] = 8'h9C;
ROM_MEM[5109] = 8'h0B;
ROM_MEM[5110] = 8'h61;
ROM_MEM[5111] = 8'h69;
ROM_MEM[5112] = 8'h65;
ROM_MEM[5113] = 8'hB6;
ROM_MEM[5114] = 8'hF0;
ROM_MEM[5115] = 8'hD6;
ROM_MEM[5116] = 8'h67;
ROM_MEM[5117] = 8'h84;
ROM_MEM[5118] = 8'h94;
ROM_MEM[5119] = 8'hD1;
ROM_MEM[5120] = 8'h26;
ROM_MEM[5121] = 8'h06;
ROM_MEM[5122] = 8'h2B;
ROM_MEM[5123] = 8'h15;
ROM_MEM[5124] = 8'h99;
ROM_MEM[5125] = 8'hB4;
ROM_MEM[5126] = 8'h9D;
ROM_MEM[5127] = 8'h9C;
ROM_MEM[5128] = 8'hB5;
ROM_MEM[5129] = 8'hB2;
ROM_MEM[5130] = 8'h79;
ROM_MEM[5131] = 8'hDA;
ROM_MEM[5132] = 8'h61;
ROM_MEM[5133] = 8'h40;
ROM_MEM[5134] = 8'hD0;
ROM_MEM[5135] = 8'hEA;
ROM_MEM[5136] = 8'h0C;
ROM_MEM[5137] = 8'h88;
ROM_MEM[5138] = 8'h4A;
ROM_MEM[5139] = 8'h3D;
ROM_MEM[5140] = 8'h89;
ROM_MEM[5141] = 8'h49;
ROM_MEM[5142] = 8'h53;
ROM_MEM[5143] = 8'h75;
ROM_MEM[5144] = 8'h87;
ROM_MEM[5145] = 8'hE2;
ROM_MEM[5146] = 8'hC1;
ROM_MEM[5147] = 8'h27;
ROM_MEM[5148] = 8'h45;
ROM_MEM[5149] = 8'hD5;
ROM_MEM[5150] = 8'h69;
ROM_MEM[5151] = 8'h8A;
ROM_MEM[5152] = 8'h07;
ROM_MEM[5153] = 8'h5B;
ROM_MEM[5154] = 8'h0D;
ROM_MEM[5155] = 8'h66;
ROM_MEM[5156] = 8'h65;
ROM_MEM[5157] = 8'h88;
ROM_MEM[5158] = 8'h4D;
ROM_MEM[5159] = 8'h8C;
ROM_MEM[5160] = 8'h2D;
ROM_MEM[5161] = 8'hE6;
ROM_MEM[5162] = 8'h66;
ROM_MEM[5163] = 8'h15;
ROM_MEM[5164] = 8'h39;
ROM_MEM[5165] = 8'hD0;
ROM_MEM[5166] = 8'h66;
ROM_MEM[5167] = 8'h96;
ROM_MEM[5168] = 8'hA9;
ROM_MEM[5169] = 8'hB9;
ROM_MEM[5170] = 8'hAD;
ROM_MEM[5171] = 8'h42;
ROM_MEM[5172] = 8'hFB;
ROM_MEM[5173] = 8'hAB;
ROM_MEM[5174] = 8'h96;
ROM_MEM[5175] = 8'hD5;
ROM_MEM[5176] = 8'h56;
ROM_MEM[5177] = 8'h17;
ROM_MEM[5178] = 8'hD3;
ROM_MEM[5179] = 8'h8C;
ROM_MEM[5180] = 8'h75;
ROM_MEM[5181] = 8'h6C;
ROM_MEM[5182] = 8'hBA;
ROM_MEM[5183] = 8'h6E;
ROM_MEM[5184] = 8'h74;
ROM_MEM[5185] = 8'h2F;
ROM_MEM[5186] = 8'hE2;
ROM_MEM[5187] = 8'h7C;
ROM_MEM[5188] = 8'h91;
ROM_MEM[5189] = 8'hA8;
ROM_MEM[5190] = 8'h31;
ROM_MEM[5191] = 8'hDD;
ROM_MEM[5192] = 8'h89;
ROM_MEM[5193] = 8'h78;
ROM_MEM[5194] = 8'h96;
ROM_MEM[5195] = 8'hED;
ROM_MEM[5196] = 8'hC2;
ROM_MEM[5197] = 8'h36;
ROM_MEM[5198] = 8'hCE;
ROM_MEM[5199] = 8'h95;
ROM_MEM[5200] = 8'h5E;
ROM_MEM[5201] = 8'h62;
ROM_MEM[5202] = 8'h1A;
ROM_MEM[5203] = 8'hDF;
ROM_MEM[5204] = 8'h1D;
ROM_MEM[5205] = 8'h78;
ROM_MEM[5206] = 8'h67;
ROM_MEM[5207] = 8'h49;
ROM_MEM[5208] = 8'h4A;
ROM_MEM[5209] = 8'h6A;
ROM_MEM[5210] = 8'hD6;
ROM_MEM[5211] = 8'hD8;
ROM_MEM[5212] = 8'hA5;
ROM_MEM[5213] = 8'h26;
ROM_MEM[5214] = 8'h39;
ROM_MEM[5215] = 8'h69;
ROM_MEM[5216] = 8'h51;
ROM_MEM[5217] = 8'h73;
ROM_MEM[5218] = 8'h36;
ROM_MEM[5219] = 8'h9B;
ROM_MEM[5220] = 8'hEC;
ROM_MEM[5221] = 8'h26;
ROM_MEM[5222] = 8'hD4;
ROM_MEM[5223] = 8'h80;
ROM_MEM[5224] = 8'h59;
ROM_MEM[5225] = 8'h35;
ROM_MEM[5226] = 8'h92;
ROM_MEM[5227] = 8'h8A;
ROM_MEM[5228] = 8'h90;
ROM_MEM[5229] = 8'h0D;
ROM_MEM[5230] = 8'hE7;
ROM_MEM[5231] = 8'h64;
ROM_MEM[5232] = 8'h8B;
ROM_MEM[5233] = 8'h72;
ROM_MEM[5234] = 8'hB2;
ROM_MEM[5235] = 8'h0E;
ROM_MEM[5236] = 8'h55;
ROM_MEM[5237] = 8'hE5;
ROM_MEM[5238] = 8'h22;
ROM_MEM[5239] = 8'hDB;
ROM_MEM[5240] = 8'h19;
ROM_MEM[5241] = 8'h4E;
ROM_MEM[5242] = 8'h7B;
ROM_MEM[5243] = 8'h64;
ROM_MEM[5244] = 8'h88;
ROM_MEM[5245] = 8'hEC;
ROM_MEM[5246] = 8'h26;
ROM_MEM[5247] = 8'hD4;
ROM_MEM[5248] = 8'h48;
ROM_MEM[5249] = 8'hE6;
ROM_MEM[5250] = 8'hBD;
ROM_MEM[5251] = 8'h96;
ROM_MEM[5252] = 8'h07;
ROM_MEM[5253] = 8'h1F;
ROM_MEM[5254] = 8'h9D;
ROM_MEM[5255] = 8'h4C;
ROM_MEM[5256] = 8'h76;
ROM_MEM[5257] = 8'hC7;
ROM_MEM[5258] = 8'h29;
ROM_MEM[5259] = 8'h82;
ROM_MEM[5260] = 8'h99;
ROM_MEM[5261] = 8'h1E;
ROM_MEM[5262] = 8'h96;
ROM_MEM[5263] = 8'h13;
ROM_MEM[5264] = 8'h3B;
ROM_MEM[5265] = 8'h09;
ROM_MEM[5266] = 8'h66;
ROM_MEM[5267] = 8'h95;
ROM_MEM[5268] = 8'hAB;
ROM_MEM[5269] = 8'h44;
ROM_MEM[5270] = 8'hDA;
ROM_MEM[5271] = 8'h20;
ROM_MEM[5272] = 8'hC9;
ROM_MEM[5273] = 8'hDB;
ROM_MEM[5274] = 8'h29;
ROM_MEM[5275] = 8'h5E;
ROM_MEM[5276] = 8'h76;
ROM_MEM[5277] = 8'h9B;
ROM_MEM[5278] = 8'hE2;
ROM_MEM[5279] = 8'hBB;
ROM_MEM[5280] = 8'h84;
ROM_MEM[5281] = 8'h4D;
ROM_MEM[5282] = 8'hD9;
ROM_MEM[5283] = 8'h6D;
ROM_MEM[5284] = 8'h5A;
ROM_MEM[5285] = 8'h2E;
ROM_MEM[5286] = 8'h1C;
ROM_MEM[5287] = 8'h9E;
ROM_MEM[5288] = 8'h25;
ROM_MEM[5289] = 8'hC7;
ROM_MEM[5290] = 8'hF9;
ROM_MEM[5291] = 8'h51;
ROM_MEM[5292] = 8'h85;
ROM_MEM[5293] = 8'h9B;
ROM_MEM[5294] = 8'h9B;
ROM_MEM[5295] = 8'hAD;
ROM_MEM[5296] = 8'h62;
ROM_MEM[5297] = 8'hE4;
ROM_MEM[5298] = 8'h28;
ROM_MEM[5299] = 8'hAA;
ROM_MEM[5300] = 8'h51;
ROM_MEM[5301] = 8'h8A;
ROM_MEM[5302] = 8'h87;
ROM_MEM[5303] = 8'h55;
ROM_MEM[5304] = 8'h9C;
ROM_MEM[5305] = 8'hBA;
ROM_MEM[5306] = 8'hED;
ROM_MEM[5307] = 8'h3A;
ROM_MEM[5308] = 8'h69;
ROM_MEM[5309] = 8'hC1;
ROM_MEM[5310] = 8'hC8;
ROM_MEM[5311] = 8'h91;
ROM_MEM[5312] = 8'h10;
ROM_MEM[5313] = 8'hE3;
ROM_MEM[5314] = 8'h38;
ROM_MEM[5315] = 8'h84;
ROM_MEM[5316] = 8'h3D;
ROM_MEM[5317] = 8'h9A;
ROM_MEM[5318] = 8'h72;
ROM_MEM[5319] = 8'h8D;
ROM_MEM[5320] = 8'hE2;
ROM_MEM[5321] = 8'h07;
ROM_MEM[5322] = 8'h22;
ROM_MEM[5323] = 8'hAA;
ROM_MEM[5324] = 8'hB6;
ROM_MEM[5325] = 8'hC3;
ROM_MEM[5326] = 8'hAD;
ROM_MEM[5327] = 8'hC9;
ROM_MEM[5328] = 8'hCF;
ROM_MEM[5329] = 8'hBC;
ROM_MEM[5330] = 8'hD2;
ROM_MEM[5331] = 8'h1C;
ROM_MEM[5332] = 8'hBF;
ROM_MEM[5333] = 8'h06;
ROM_MEM[5334] = 8'hAF;
ROM_MEM[5335] = 8'hD0;
ROM_MEM[5336] = 8'h49;
ROM_MEM[5337] = 8'hB2;
ROM_MEM[5338] = 8'h82;
ROM_MEM[5339] = 8'h3E;
ROM_MEM[5340] = 8'h65;
ROM_MEM[5341] = 8'hD2;
ROM_MEM[5342] = 8'hA4;
ROM_MEM[5343] = 8'hAA;
ROM_MEM[5344] = 8'h01;
ROM_MEM[5345] = 8'h6A;
ROM_MEM[5346] = 8'h95;
ROM_MEM[5347] = 8'h72;
ROM_MEM[5348] = 8'h40;
ROM_MEM[5349] = 8'hAE;
ROM_MEM[5350] = 8'hD6;
ROM_MEM[5351] = 8'h43;
ROM_MEM[5352] = 8'hAB;
ROM_MEM[5353] = 8'h2E;
ROM_MEM[5354] = 8'hFA;
ROM_MEM[5355] = 8'hD4;
ROM_MEM[5356] = 8'h93;
ROM_MEM[5357] = 8'h2E;
ROM_MEM[5358] = 8'h35;
ROM_MEM[5359] = 8'h07;
ROM_MEM[5360] = 8'h5B;
ROM_MEM[5361] = 8'hD3;
ROM_MEM[5362] = 8'h4C;
ROM_MEM[5363] = 8'hB6;
ROM_MEM[5364] = 8'hE4;
ROM_MEM[5365] = 8'h34;
ROM_MEM[5366] = 8'h72;
ROM_MEM[5367] = 8'h54;
ROM_MEM[5368] = 8'hA7;
ROM_MEM[5369] = 8'hCD;
ROM_MEM[5370] = 8'h91;
ROM_MEM[5371] = 8'h52;
ROM_MEM[5372] = 8'hEE;
ROM_MEM[5373] = 8'h4A;
ROM_MEM[5374] = 8'hA9;
ROM_MEM[5375] = 8'hB9;
ROM_MEM[5376] = 8'h47;
ROM_MEM[5377] = 8'hAA;
ROM_MEM[5378] = 8'hC1;
ROM_MEM[5379] = 8'h56;
ROM_MEM[5380] = 8'hB5;
ROM_MEM[5381] = 8'hD2;
ROM_MEM[5382] = 8'h2E;
ROM_MEM[5383] = 8'hB9;
ROM_MEM[5384] = 8'hF8;
ROM_MEM[5385] = 8'hAC;
ROM_MEM[5386] = 8'hB6;
ROM_MEM[5387] = 8'h4C;
ROM_MEM[5388] = 8'h12;
ROM_MEM[5389] = 8'h80;
ROM_MEM[5390] = 8'h66;
ROM_MEM[5391] = 8'hCA;
ROM_MEM[5392] = 8'h04;
ROM_MEM[5393] = 8'h90;
ROM_MEM[5394] = 8'hD4;
ROM_MEM[5395] = 8'h9A;
ROM_MEM[5396] = 8'h01;
ROM_MEM[5397] = 8'hA6;
ROM_MEM[5398] = 8'h75;
ROM_MEM[5399] = 8'h3E;
ROM_MEM[5400] = 8'h52;
ROM_MEM[5401] = 8'hC9;
ROM_MEM[5402] = 8'h91;
ROM_MEM[5403] = 8'h65;
ROM_MEM[5404] = 8'h16;
ROM_MEM[5405] = 8'hF6;
ROM_MEM[5406] = 8'hA8;
ROM_MEM[5407] = 8'hA5;
ROM_MEM[5408] = 8'h79;
ROM_MEM[5409] = 8'h74;
ROM_MEM[5410] = 8'hB1;
ROM_MEM[5411] = 8'hBB;
ROM_MEM[5412] = 8'hA3;
ROM_MEM[5413] = 8'h95;
ROM_MEM[5414] = 8'hE9;
ROM_MEM[5415] = 8'hBE;
ROM_MEM[5416] = 8'h49;
ROM_MEM[5417] = 8'hCD;
ROM_MEM[5418] = 8'h96;
ROM_MEM[5419] = 8'h9E;
ROM_MEM[5420] = 8'h4F;
ROM_MEM[5421] = 8'hDA;
ROM_MEM[5422] = 8'h84;
ROM_MEM[5423] = 8'hB4;
ROM_MEM[5424] = 8'h1D;
ROM_MEM[5425] = 8'h6A;
ROM_MEM[5426] = 8'h7D;
ROM_MEM[5427] = 8'h11;
ROM_MEM[5428] = 8'h19;
ROM_MEM[5429] = 8'h16;
ROM_MEM[5430] = 8'h17;
ROM_MEM[5431] = 8'hA0;
ROM_MEM[5432] = 8'h00;
ROM_MEM[5433] = 8'hA3;
ROM_MEM[5434] = 8'hB5;
ROM_MEM[5435] = 8'h1F;
ROM_MEM[5436] = 8'hBE;
ROM_MEM[5437] = 8'hF7;
ROM_MEM[5438] = 8'hC9;
ROM_MEM[5439] = 8'h31;
ROM_MEM[5440] = 8'h4E;
ROM_MEM[5441] = 8'h72;
ROM_MEM[5442] = 8'h98;
ROM_MEM[5443] = 8'hB6;
ROM_MEM[5444] = 8'hA6;
ROM_MEM[5445] = 8'h57;
ROM_MEM[5446] = 8'h69;
ROM_MEM[5447] = 8'hCA;
ROM_MEM[5448] = 8'h62;
ROM_MEM[5449] = 8'h46;
ROM_MEM[5450] = 8'hCF;
ROM_MEM[5451] = 8'h28;
ROM_MEM[5452] = 8'hD6;
ROM_MEM[5453] = 8'h3A;
ROM_MEM[5454] = 8'h8D;
ROM_MEM[5455] = 8'h19;
ROM_MEM[5456] = 8'h4D;
ROM_MEM[5457] = 8'hB3;
ROM_MEM[5458] = 8'h45;
ROM_MEM[5459] = 8'hEB;
ROM_MEM[5460] = 8'h0E;
ROM_MEM[5461] = 8'hAE;
ROM_MEM[5462] = 8'h06;
ROM_MEM[5463] = 8'hEF;
ROM_MEM[5464] = 8'h31;
ROM_MEM[5465] = 8'h4A;
ROM_MEM[5466] = 8'h5A;
ROM_MEM[5467] = 8'hA4;
ROM_MEM[5468] = 8'hEC;
ROM_MEM[5469] = 8'hAB;
ROM_MEM[5470] = 8'h93;
ROM_MEM[5471] = 8'hA5;
ROM_MEM[5472] = 8'h71;
ROM_MEM[5473] = 8'hF2;
ROM_MEM[5474] = 8'h52;
ROM_MEM[5475] = 8'hC8;
ROM_MEM[5476] = 8'h75;
ROM_MEM[5477] = 8'hD6;
ROM_MEM[5478] = 8'hA8;
ROM_MEM[5479] = 8'h0C;
ROM_MEM[5480] = 8'hF0;
ROM_MEM[5481] = 8'hB5;
ROM_MEM[5482] = 8'h82;
ROM_MEM[5483] = 8'h01;
ROM_MEM[5484] = 8'hBE;
ROM_MEM[5485] = 8'h4C;
ROM_MEM[5486] = 8'h12;
ROM_MEM[5487] = 8'h20;
ROM_MEM[5488] = 8'hB8;
ROM_MEM[5489] = 8'h0C;
ROM_MEM[5490] = 8'h02;
ROM_MEM[5491] = 8'h04;
ROM_MEM[5492] = 8'h13;
ROM_MEM[5493] = 8'h8A;
ROM_MEM[5494] = 8'h80;
ROM_MEM[5495] = 8'h80;
ROM_MEM[5496] = 8'h44;
ROM_MEM[5497] = 8'h1E;
ROM_MEM[5498] = 8'hE0;
ROM_MEM[5499] = 8'hCB;
ROM_MEM[5500] = 8'h24;
ROM_MEM[5501] = 8'h89;
ROM_MEM[5502] = 8'h6A;
ROM_MEM[5503] = 8'hE4;
ROM_MEM[5504] = 8'h3C;
ROM_MEM[5505] = 8'hCD;
ROM_MEM[5506] = 8'hDD;
ROM_MEM[5507] = 8'h04;
ROM_MEM[5508] = 8'hA5;
ROM_MEM[5509] = 8'h48;
ROM_MEM[5510] = 8'hF7;
ROM_MEM[5511] = 8'h10;
ROM_MEM[5512] = 8'hA7;
ROM_MEM[5513] = 8'h13;
ROM_MEM[5514] = 8'h98;
ROM_MEM[5515] = 8'h50;
ROM_MEM[5516] = 8'hDC;
ROM_MEM[5517] = 8'h2D;
ROM_MEM[5518] = 8'h44;
ROM_MEM[5519] = 8'h69;
ROM_MEM[5520] = 8'h22;
ROM_MEM[5521] = 8'h43;
ROM_MEM[5522] = 8'h67;
ROM_MEM[5523] = 8'hF5;
ROM_MEM[5524] = 8'h34;
ROM_MEM[5525] = 8'hA7;
ROM_MEM[5526] = 8'h03;
ROM_MEM[5527] = 8'h4B;
ROM_MEM[5528] = 8'hEB;
ROM_MEM[5529] = 8'hC2;
ROM_MEM[5530] = 8'h4C;
ROM_MEM[5531] = 8'h94;
ROM_MEM[5532] = 8'h0E;
ROM_MEM[5533] = 8'hAC;
ROM_MEM[5534] = 8'hAE;
ROM_MEM[5535] = 8'h28;
ROM_MEM[5536] = 8'h6F;
ROM_MEM[5537] = 8'hAD;
ROM_MEM[5538] = 8'hBD;
ROM_MEM[5539] = 8'hD0;
ROM_MEM[5540] = 8'h95;
ROM_MEM[5541] = 8'hBA;
ROM_MEM[5542] = 8'hB9;
ROM_MEM[5543] = 8'hB4;
ROM_MEM[5544] = 8'hCA;
ROM_MEM[5545] = 8'h42;
ROM_MEM[5546] = 8'h57;
ROM_MEM[5547] = 8'h1A;
ROM_MEM[5548] = 8'h77;
ROM_MEM[5549] = 8'h0A;
ROM_MEM[5550] = 8'hCB;
ROM_MEM[5551] = 8'h0B;
ROM_MEM[5552] = 8'h9F;
ROM_MEM[5553] = 8'h31;
ROM_MEM[5554] = 8'hD0;
ROM_MEM[5555] = 8'h2C;
ROM_MEM[5556] = 8'hEB;
ROM_MEM[5557] = 8'h16;
ROM_MEM[5558] = 8'h6A;
ROM_MEM[5559] = 8'h45;
ROM_MEM[5560] = 8'h47;
ROM_MEM[5561] = 8'h0D;
ROM_MEM[5562] = 8'hAD;
ROM_MEM[5563] = 8'h13;
ROM_MEM[5564] = 8'hA4;
ROM_MEM[5565] = 8'h69;
ROM_MEM[5566] = 8'h15;
ROM_MEM[5567] = 8'hDD;
ROM_MEM[5568] = 8'hAD;
ROM_MEM[5569] = 8'h8E;
ROM_MEM[5570] = 8'hD3;
ROM_MEM[5571] = 8'h67;
ROM_MEM[5572] = 8'h4C;
ROM_MEM[5573] = 8'h35;
ROM_MEM[5574] = 8'h36;
ROM_MEM[5575] = 8'h29;
ROM_MEM[5576] = 8'h0E;
ROM_MEM[5577] = 8'h28;
ROM_MEM[5578] = 8'h50;
ROM_MEM[5579] = 8'h34;
ROM_MEM[5580] = 8'h00;
ROM_MEM[5581] = 8'h93;
ROM_MEM[5582] = 8'h12;
ROM_MEM[5583] = 8'h27;
ROM_MEM[5584] = 8'h60;
ROM_MEM[5585] = 8'h4A;
ROM_MEM[5586] = 8'hA5;
ROM_MEM[5587] = 8'h41;
ROM_MEM[5588] = 8'h76;
ROM_MEM[5589] = 8'h95;
ROM_MEM[5590] = 8'h2A;
ROM_MEM[5591] = 8'h9A;
ROM_MEM[5592] = 8'hB1;
ROM_MEM[5593] = 8'h0F;
ROM_MEM[5594] = 8'h51;
ROM_MEM[5595] = 8'h7D;
ROM_MEM[5596] = 8'h86;
ROM_MEM[5597] = 8'hB4;
ROM_MEM[5598] = 8'hA7;
ROM_MEM[5599] = 8'h59;
ROM_MEM[5600] = 8'h44;
ROM_MEM[5601] = 8'h4D;
ROM_MEM[5602] = 8'hE9;
ROM_MEM[5603] = 8'h19;
ROM_MEM[5604] = 8'h96;
ROM_MEM[5605] = 8'h76;
ROM_MEM[5606] = 8'h51;
ROM_MEM[5607] = 8'hC5;
ROM_MEM[5608] = 8'h77;
ROM_MEM[5609] = 8'h56;
ROM_MEM[5610] = 8'hD5;
ROM_MEM[5611] = 8'h92;
ROM_MEM[5612] = 8'h41;
ROM_MEM[5613] = 8'h97;
ROM_MEM[5614] = 8'h94;
ROM_MEM[5615] = 8'hE5;
ROM_MEM[5616] = 8'h9D;
ROM_MEM[5617] = 8'h6B;
ROM_MEM[5618] = 8'h06;
ROM_MEM[5619] = 8'hDB;
ROM_MEM[5620] = 8'h62;
ROM_MEM[5621] = 8'h66;
ROM_MEM[5622] = 8'h66;
ROM_MEM[5623] = 8'hD4;
ROM_MEM[5624] = 8'h6D;
ROM_MEM[5625] = 8'h5C;
ROM_MEM[5626] = 8'hEB;
ROM_MEM[5627] = 8'h15;
ROM_MEM[5628] = 8'h6A;
ROM_MEM[5629] = 8'h51;
ROM_MEM[5630] = 8'hDB;
ROM_MEM[5631] = 8'h71;
ROM_MEM[5632] = 8'h2D;
ROM_MEM[5633] = 8'h57;
ROM_MEM[5634] = 8'h98;
ROM_MEM[5635] = 8'h69;
ROM_MEM[5636] = 8'h69;
ROM_MEM[5637] = 8'h06;
ROM_MEM[5638] = 8'h60;
ROM_MEM[5639] = 8'hA1;
ROM_MEM[5640] = 8'h86;
ROM_MEM[5641] = 8'h00;
ROM_MEM[5642] = 8'hA4;
ROM_MEM[5643] = 8'h44;
ROM_MEM[5644] = 8'h41;
ROM_MEM[5645] = 8'h01;
ROM_MEM[5646] = 8'h09;
ROM_MEM[5647] = 8'hB2;
ROM_MEM[5648] = 8'h14;
ROM_MEM[5649] = 8'h71;
ROM_MEM[5650] = 8'h87;
ROM_MEM[5651] = 8'hF2;
ROM_MEM[5652] = 8'h34;
ROM_MEM[5653] = 8'h8F;
ROM_MEM[5654] = 8'hB2;
ROM_MEM[5655] = 8'hA8;
ROM_MEM[5656] = 8'hE1;
ROM_MEM[5657] = 8'hD5;
ROM_MEM[5658] = 8'h20;
ROM_MEM[5659] = 8'h33;
ROM_MEM[5660] = 8'hC9;
ROM_MEM[5661] = 8'hA1;
ROM_MEM[5662] = 8'h46;
ROM_MEM[5663] = 8'h35;
ROM_MEM[5664] = 8'h15;
ROM_MEM[5665] = 8'h4F;
ROM_MEM[5666] = 8'hC7;
ROM_MEM[5667] = 8'h83;
ROM_MEM[5668] = 8'h69;
ROM_MEM[5669] = 8'h5E;
ROM_MEM[5670] = 8'hC2;
ROM_MEM[5671] = 8'hBA;
ROM_MEM[5672] = 8'h93;
ROM_MEM[5673] = 8'h0E;
ROM_MEM[5674] = 8'hB6;
ROM_MEM[5675] = 8'h45;
ROM_MEM[5676] = 8'h0D;
ROM_MEM[5677] = 8'hB1;
ROM_MEM[5678] = 8'h4B;
ROM_MEM[5679] = 8'h12;
ROM_MEM[5680] = 8'hA4;
ROM_MEM[5681] = 8'h16;
ROM_MEM[5682] = 8'h34;
ROM_MEM[5683] = 8'hC8;
ROM_MEM[5684] = 8'h2A;
ROM_MEM[5685] = 8'h56;
ROM_MEM[5686] = 8'h50;
ROM_MEM[5687] = 8'hAA;
ROM_MEM[5688] = 8'h13;
ROM_MEM[5689] = 8'h55;
ROM_MEM[5690] = 8'h2B;
ROM_MEM[5691] = 8'hCB;
ROM_MEM[5692] = 8'h41;
ROM_MEM[5693] = 8'hAE;
ROM_MEM[5694] = 8'hD6;
ROM_MEM[5695] = 8'h54;
ROM_MEM[5696] = 8'h25;
ROM_MEM[5697] = 8'h13;
ROM_MEM[5698] = 8'h2D;
ROM_MEM[5699] = 8'h26;
ROM_MEM[5700] = 8'h39;
ROM_MEM[5701] = 8'hB3;
ROM_MEM[5702] = 8'h9E;
ROM_MEM[5703] = 8'h49;
ROM_MEM[5704] = 8'h72;
ROM_MEM[5705] = 8'h98;
ROM_MEM[5706] = 8'h96;
ROM_MEM[5707] = 8'hD3;
ROM_MEM[5708] = 8'hB4;
ROM_MEM[5709] = 8'h2A;
ROM_MEM[5710] = 8'hEA;
ROM_MEM[5711] = 8'h61;
ROM_MEM[5712] = 8'h9A;
ROM_MEM[5713] = 8'h1B;
ROM_MEM[5714] = 8'hF7;
ROM_MEM[5715] = 8'hB2;
ROM_MEM[5716] = 8'hA6;
ROM_MEM[5717] = 8'h8B;
ROM_MEM[5718] = 8'h2D;
ROM_MEM[5719] = 8'h76;
ROM_MEM[5720] = 8'hD3;
ROM_MEM[5721] = 8'h92;
ROM_MEM[5722] = 8'hD3;
ROM_MEM[5723] = 8'h26;
ROM_MEM[5724] = 8'h2E;
ROM_MEM[5725] = 8'hD9;
ROM_MEM[5726] = 8'h8C;
ROM_MEM[5727] = 8'h08;
ROM_MEM[5728] = 8'h6B;
ROM_MEM[5729] = 8'hE2;
ROM_MEM[5730] = 8'h84;
ROM_MEM[5731] = 8'hA6;
ROM_MEM[5732] = 8'hCC;
ROM_MEM[5733] = 8'hB2;
ROM_MEM[5734] = 8'hB4;
ROM_MEM[5735] = 8'h75;
ROM_MEM[5736] = 8'h62;
ROM_MEM[5737] = 8'h2B;
ROM_MEM[5738] = 8'hF7;
ROM_MEM[5739] = 8'h75;
ROM_MEM[5740] = 8'hE7;
ROM_MEM[5741] = 8'h36;
ROM_MEM[5742] = 8'h8D;
ROM_MEM[5743] = 8'hCD;
ROM_MEM[5744] = 8'h66;
ROM_MEM[5745] = 8'h93;
ROM_MEM[5746] = 8'hDC;
ROM_MEM[5747] = 8'hDE;
ROM_MEM[5748] = 8'h34;
ROM_MEM[5749] = 8'hBE;
ROM_MEM[5750] = 8'h8B;
ROM_MEM[5751] = 8'h76;
ROM_MEM[5752] = 8'h67;
ROM_MEM[5753] = 8'h6D;
ROM_MEM[5754] = 8'h5C;
ROM_MEM[5755] = 8'hF4;
ROM_MEM[5756] = 8'h6B;
ROM_MEM[5757] = 8'h4D;
ROM_MEM[5758] = 8'hDC;
ROM_MEM[5759] = 8'hCD;
ROM_MEM[5760] = 8'h76;
ROM_MEM[5761] = 8'h93;
ROM_MEM[5762] = 8'h0A;
ROM_MEM[5763] = 8'h77;
ROM_MEM[5764] = 8'h8B;
ROM_MEM[5765] = 8'h64;
ROM_MEM[5766] = 8'hCF;
ROM_MEM[5767] = 8'h85;
ROM_MEM[5768] = 8'hCF;
ROM_MEM[5769] = 8'h9A;
ROM_MEM[5770] = 8'h6A;
ROM_MEM[5771] = 8'h52;
ROM_MEM[5772] = 8'h65;
ROM_MEM[5773] = 8'h37;
ROM_MEM[5774] = 8'h36;
ROM_MEM[5775] = 8'h29;
ROM_MEM[5776] = 8'h9D;
ROM_MEM[5777] = 8'hEE;
ROM_MEM[5778] = 8'h0C;
ROM_MEM[5779] = 8'hD3;
ROM_MEM[5780] = 8'hE8;
ROM_MEM[5781] = 8'h28;
ROM_MEM[5782] = 8'h6B;
ROM_MEM[5783] = 8'hBA;
ROM_MEM[5784] = 8'h54;
ROM_MEM[5785] = 8'hEA;
ROM_MEM[5786] = 8'hA0;
ROM_MEM[5787] = 8'h93;
ROM_MEM[5788] = 8'hEF;
ROM_MEM[5789] = 8'h09;
ROM_MEM[5790] = 8'hA7;
ROM_MEM[5791] = 8'hA4;
ROM_MEM[5792] = 8'h83;
ROM_MEM[5793] = 8'hCA;
ROM_MEM[5794] = 8'h6D;
ROM_MEM[5795] = 8'h92;
ROM_MEM[5796] = 8'h53;
ROM_MEM[5797] = 8'h17;
ROM_MEM[5798] = 8'h37;
ROM_MEM[5799] = 8'hBA;
ROM_MEM[5800] = 8'h26;
ROM_MEM[5801] = 8'h19;
ROM_MEM[5802] = 8'h71;
ROM_MEM[5803] = 8'hF7;
ROM_MEM[5804] = 8'hB2;
ROM_MEM[5805] = 8'hA8;
ROM_MEM[5806] = 8'h16;
ROM_MEM[5807] = 8'hB5;
ROM_MEM[5808] = 8'h34;
ROM_MEM[5809] = 8'hBC;
ROM_MEM[5810] = 8'hE9;
ROM_MEM[5811] = 8'hA2;
ROM_MEM[5812] = 8'h6B;
ROM_MEM[5813] = 8'hB1;
ROM_MEM[5814] = 8'h94;
ROM_MEM[5815] = 8'hD4;
ROM_MEM[5816] = 8'h25;
ROM_MEM[5817] = 8'h8D;
ROM_MEM[5818] = 8'hAE;
ROM_MEM[5819] = 8'h35;
ROM_MEM[5820] = 8'h82;
ROM_MEM[5821] = 8'h5C;
ROM_MEM[5822] = 8'hEA;
ROM_MEM[5823] = 8'h14;
ROM_MEM[5824] = 8'hA6;
ROM_MEM[5825] = 8'h5B;
ROM_MEM[5826] = 8'h4C;
ROM_MEM[5827] = 8'h49;
ROM_MEM[5828] = 8'h6B;
ROM_MEM[5829] = 8'h75;
ROM_MEM[5830] = 8'h98;
ROM_MEM[5831] = 8'h1E;
ROM_MEM[5832] = 8'h35;
ROM_MEM[5833] = 8'h29;
ROM_MEM[5834] = 8'hD3;
ROM_MEM[5835] = 8'hCB;
ROM_MEM[5836] = 8'h62;
ROM_MEM[5837] = 8'hBB;
ROM_MEM[5838] = 8'h71;
ROM_MEM[5839] = 8'h97;
ROM_MEM[5840] = 8'h89;
ROM_MEM[5841] = 8'h39;
ROM_MEM[5842] = 8'h85;
ROM_MEM[5843] = 8'h2B;
ROM_MEM[5844] = 8'hDA;
ROM_MEM[5845] = 8'hDD;
ROM_MEM[5846] = 8'h9A;
ROM_MEM[5847] = 8'h93;
ROM_MEM[5848] = 8'h26;
ROM_MEM[5849] = 8'hBE;
ROM_MEM[5850] = 8'h58;
ROM_MEM[5851] = 8'hF6;
ROM_MEM[5852] = 8'h0C;
ROM_MEM[5853] = 8'hAD;
ROM_MEM[5854] = 8'h9D;
ROM_MEM[5855] = 8'hF8;
ROM_MEM[5856] = 8'h16;
ROM_MEM[5857] = 8'h49;
ROM_MEM[5858] = 8'hB2;
ROM_MEM[5859] = 8'hA9;
ROM_MEM[5860] = 8'hE1;
ROM_MEM[5861] = 8'hE2;
ROM_MEM[5862] = 8'h86;
ROM_MEM[5863] = 8'hB4;
ROM_MEM[5864] = 8'h90;
ROM_MEM[5865] = 8'hF6;
ROM_MEM[5866] = 8'hA5;
ROM_MEM[5867] = 8'h8B;
ROM_MEM[5868] = 8'hAB;
ROM_MEM[5869] = 8'h26;
ROM_MEM[5870] = 8'h4C;
ROM_MEM[5871] = 8'h3A;
ROM_MEM[5872] = 8'hE7;
ROM_MEM[5873] = 8'h2C;
ROM_MEM[5874] = 8'hBE;
ROM_MEM[5875] = 8'h29;
ROM_MEM[5876] = 8'h2B;
ROM_MEM[5877] = 8'h75;
ROM_MEM[5878] = 8'h9F;
ROM_MEM[5879] = 8'h37;
ROM_MEM[5880] = 8'h84;
ROM_MEM[5881] = 8'h66;
ROM_MEM[5882] = 8'hB4;
ROM_MEM[5883] = 8'h55;
ROM_MEM[5884] = 8'hFC;
ROM_MEM[5885] = 8'hCE;
ROM_MEM[5886] = 8'h12;
ROM_MEM[5887] = 8'hAB;
ROM_MEM[5888] = 8'hF6;
ROM_MEM[5889] = 8'hE0;
ROM_MEM[5890] = 8'h8C;
ROM_MEM[5891] = 8'h27;
ROM_MEM[5892] = 8'h43;
ROM_MEM[5893] = 8'hE9;
ROM_MEM[5894] = 8'h56;
ROM_MEM[5895] = 8'h4C;
ROM_MEM[5896] = 8'h33;
ROM_MEM[5897] = 8'hE6;
ROM_MEM[5898] = 8'h36;
ROM_MEM[5899] = 8'h65;
ROM_MEM[5900] = 8'h66;
ROM_MEM[5901] = 8'h77;
ROM_MEM[5902] = 8'h32;
ROM_MEM[5903] = 8'h1D;
ROM_MEM[5904] = 8'hDD;
ROM_MEM[5905] = 8'hB4;
ROM_MEM[5906] = 8'h11;
ROM_MEM[5907] = 8'h55;
ROM_MEM[5908] = 8'hA9;
ROM_MEM[5909] = 8'hB2;
ROM_MEM[5910] = 8'hF2;
ROM_MEM[5911] = 8'hB2;
ROM_MEM[5912] = 8'h7A;
ROM_MEM[5913] = 8'h12;
ROM_MEM[5914] = 8'hE5;
ROM_MEM[5915] = 8'hCC;
ROM_MEM[5916] = 8'hBA;
ROM_MEM[5917] = 8'hCB;
ROM_MEM[5918] = 8'h6D;
ROM_MEM[5919] = 8'h49;
ROM_MEM[5920] = 8'hCC;
ROM_MEM[5921] = 8'h32;
ROM_MEM[5922] = 8'h6B;
ROM_MEM[5923] = 8'h8F;
ROM_MEM[5924] = 8'hA0;
ROM_MEM[5925] = 8'h44;
ROM_MEM[5926] = 8'h8E;
ROM_MEM[5927] = 8'h88;
ROM_MEM[5928] = 8'h8A;
ROM_MEM[5929] = 8'h5D;
ROM_MEM[5930] = 8'hC2;
ROM_MEM[5931] = 8'h1C;
ROM_MEM[5932] = 8'hC5;
ROM_MEM[5933] = 8'h52;
ROM_MEM[5934] = 8'hBB;
ROM_MEM[5935] = 8'h76;
ROM_MEM[5936] = 8'h88;
ROM_MEM[5937] = 8'h8A;
ROM_MEM[5938] = 8'h23;
ROM_MEM[5939] = 8'h0F;
ROM_MEM[5940] = 8'h8F;
ROM_MEM[5941] = 8'h34;
ROM_MEM[5942] = 8'h21;
ROM_MEM[5943] = 8'hAA;
ROM_MEM[5944] = 8'h9E;
ROM_MEM[5945] = 8'hDC;
ROM_MEM[5946] = 8'hDC;
ROM_MEM[5947] = 8'h9D;
ROM_MEM[5948] = 8'hB9;
ROM_MEM[5949] = 8'h28;
ROM_MEM[5950] = 8'h09;
ROM_MEM[5951] = 8'h8D;
ROM_MEM[5952] = 8'h8C;
ROM_MEM[5953] = 8'h8C;
ROM_MEM[5954] = 8'hF5;
ROM_MEM[5955] = 8'h00;
ROM_MEM[5956] = 8'hA5;
ROM_MEM[5957] = 8'h3A;
ROM_MEM[5958] = 8'h51;
ROM_MEM[5959] = 8'hC3;
ROM_MEM[5960] = 8'h4D;
ROM_MEM[5961] = 8'hC1;
ROM_MEM[5962] = 8'h6A;
ROM_MEM[5963] = 8'hBC;
ROM_MEM[5964] = 8'h98;
ROM_MEM[5965] = 8'h24;
ROM_MEM[5966] = 8'h2F;
ROM_MEM[5967] = 8'h49;
ROM_MEM[5968] = 8'hD7;
ROM_MEM[5969] = 8'hB5;
ROM_MEM[5970] = 8'h94;
ROM_MEM[5971] = 8'h02;
ROM_MEM[5972] = 8'h10;
ROM_MEM[5973] = 8'h80;
ROM_MEM[5974] = 8'h66;
ROM_MEM[5975] = 8'hD5;
ROM_MEM[5976] = 8'h06;
ROM_MEM[5977] = 8'h93;
ROM_MEM[5978] = 8'h0C;
ROM_MEM[5979] = 8'hB7;
ROM_MEM[5980] = 8'h99;
ROM_MEM[5981] = 8'h2B;
ROM_MEM[5982] = 8'h3E;
ROM_MEM[5983] = 8'h64;
ROM_MEM[5984] = 8'h8D;
ROM_MEM[5985] = 8'hD4;
ROM_MEM[5986] = 8'h56;
ROM_MEM[5987] = 8'h61;
ROM_MEM[5988] = 8'h6B;
ROM_MEM[5989] = 8'h91;
ROM_MEM[5990] = 8'h3D;
ROM_MEM[5991] = 8'h52;
ROM_MEM[5992] = 8'hA5;
ROM_MEM[5993] = 8'h67;
ROM_MEM[5994] = 8'hA2;
ROM_MEM[5995] = 8'h43;
ROM_MEM[5996] = 8'h34;
ROM_MEM[5997] = 8'hA7;
ROM_MEM[5998] = 8'hE9;
ROM_MEM[5999] = 8'h39;
ROM_MEM[6000] = 8'h09;
ROM_MEM[6001] = 8'h0F;
ROM_MEM[6002] = 8'h5E;
ROM_MEM[6003] = 8'h9D;
ROM_MEM[6004] = 8'hA6;
ROM_MEM[6005] = 8'h4F;
ROM_MEM[6006] = 8'h39;
ROM_MEM[6007] = 8'h3C;
ROM_MEM[6008] = 8'h78;
ROM_MEM[6009] = 8'h0D;
ROM_MEM[6010] = 8'h9A;
ROM_MEM[6011] = 8'hB6;
ROM_MEM[6012] = 8'h65;
ROM_MEM[6013] = 8'hB9;
ROM_MEM[6014] = 8'h91;
ROM_MEM[6015] = 8'h35;
ROM_MEM[6016] = 8'h52;
ROM_MEM[6017] = 8'h70;
ROM_MEM[6018] = 8'hBB;
ROM_MEM[6019] = 8'h2D;
ROM_MEM[6020] = 8'h25;
ROM_MEM[6021] = 8'h78;
ROM_MEM[6022] = 8'hE1;
ROM_MEM[6023] = 8'h15;
ROM_MEM[6024] = 8'h91;
ROM_MEM[6025] = 8'hB4;
ROM_MEM[6026] = 8'h8D;
ROM_MEM[6027] = 8'h3D;
ROM_MEM[6028] = 8'h95;
ROM_MEM[6029] = 8'h49;
ROM_MEM[6030] = 8'hA8;
ROM_MEM[6031] = 8'h38;
ROM_MEM[6032] = 8'h71;
ROM_MEM[6033] = 8'h40;
ROM_MEM[6034] = 8'hA3;
ROM_MEM[6035] = 8'h1E;
ROM_MEM[6036] = 8'h0E;
ROM_MEM[6037] = 8'h18;
ROM_MEM[6038] = 8'h44;
ROM_MEM[6039] = 8'hD8;
ROM_MEM[6040] = 8'h01;
ROM_MEM[6041] = 8'h83;
ROM_MEM[6042] = 8'h8B;
ROM_MEM[6043] = 8'h16;
ROM_MEM[6044] = 8'hAA;
ROM_MEM[6045] = 8'h4B;
ROM_MEM[6046] = 8'h91;
ROM_MEM[6047] = 8'h14;
ROM_MEM[6048] = 8'h6F;
ROM_MEM[6049] = 8'hBB;
ROM_MEM[6050] = 8'hF0;
ROM_MEM[6051] = 8'h1C;
ROM_MEM[6052] = 8'hD0;
ROM_MEM[6053] = 8'hDB;
ROM_MEM[6054] = 8'hCA;
ROM_MEM[6055] = 8'hED;
ROM_MEM[6056] = 8'hC1;
ROM_MEM[6057] = 8'h53;
ROM_MEM[6058] = 8'h70;
ROM_MEM[6059] = 8'hBB;
ROM_MEM[6060] = 8'h6C;
ROM_MEM[6061] = 8'hA9;
ROM_MEM[6062] = 8'h07;
ROM_MEM[6063] = 8'hCB;
ROM_MEM[6064] = 8'h51;
ROM_MEM[6065] = 8'h73;
ROM_MEM[6066] = 8'h73;
ROM_MEM[6067] = 8'hDC;
ROM_MEM[6068] = 8'h1D;
ROM_MEM[6069] = 8'hB4;
ROM_MEM[6070] = 8'h04;
ROM_MEM[6071] = 8'hED;
ROM_MEM[6072] = 8'hE8;
ROM_MEM[6073] = 8'h4E;
ROM_MEM[6074] = 8'hBD;
ROM_MEM[6075] = 8'hD0;
ROM_MEM[6076] = 8'hE2;
ROM_MEM[6077] = 8'h64;
ROM_MEM[6078] = 8'h27;
ROM_MEM[6079] = 8'hD7;
ROM_MEM[6080] = 8'hCE;
ROM_MEM[6081] = 8'h42;
ROM_MEM[6082] = 8'hE6;
ROM_MEM[6083] = 8'h24;
ROM_MEM[6084] = 8'h1F;
ROM_MEM[6085] = 8'h0F;
ROM_MEM[6086] = 8'h9B;
ROM_MEM[6087] = 8'h03;
ROM_MEM[6088] = 8'h1D;
ROM_MEM[6089] = 8'h19;
ROM_MEM[6090] = 8'hB5;
ROM_MEM[6091] = 8'h32;
ROM_MEM[6092] = 8'h33;
ROM_MEM[6093] = 8'h05;
ROM_MEM[6094] = 8'hB2;
ROM_MEM[6095] = 8'h08;
ROM_MEM[6096] = 8'hAE;
ROM_MEM[6097] = 8'hF2;
ROM_MEM[6098] = 8'hB4;
ROM_MEM[6099] = 8'h6C;
ROM_MEM[6100] = 8'hC4;
ROM_MEM[6101] = 8'hCC;
ROM_MEM[6102] = 8'hD4;
ROM_MEM[6103] = 8'hDB;
ROM_MEM[6104] = 8'hC3;
ROM_MEM[6105] = 8'h16;
ROM_MEM[6106] = 8'h03;
ROM_MEM[6107] = 8'h22;
ROM_MEM[6108] = 8'h75;
ROM_MEM[6109] = 8'h4D;
ROM_MEM[6110] = 8'h5C;
ROM_MEM[6111] = 8'h92;
ROM_MEM[6112] = 8'h9C;
ROM_MEM[6113] = 8'h99;
ROM_MEM[6114] = 8'h29;
ROM_MEM[6115] = 8'hAB;
ROM_MEM[6116] = 8'h89;
ROM_MEM[6117] = 8'hD9;
ROM_MEM[6118] = 8'h51;
ROM_MEM[6119] = 8'hC5;
ROM_MEM[6120] = 8'hB4;
ROM_MEM[6121] = 8'hE2;
ROM_MEM[6122] = 8'h66;
ROM_MEM[6123] = 8'hD5;
ROM_MEM[6124] = 8'hC6;
ROM_MEM[6125] = 8'hA6;
ROM_MEM[6126] = 8'hB9;
ROM_MEM[6127] = 8'h8A;
ROM_MEM[6128] = 8'h8B;
ROM_MEM[6129] = 8'h9F;
ROM_MEM[6130] = 8'h02;
ROM_MEM[6131] = 8'hA5;
ROM_MEM[6132] = 8'h5F;
ROM_MEM[6133] = 8'h3B;
ROM_MEM[6134] = 8'h71;
ROM_MEM[6135] = 8'h71;
ROM_MEM[6136] = 8'h54;
ROM_MEM[6137] = 8'h66;
ROM_MEM[6138] = 8'hE6;
ROM_MEM[6139] = 8'h95;
ROM_MEM[6140] = 8'hDA;
ROM_MEM[6141] = 8'h64;
ROM_MEM[6142] = 8'h99;
ROM_MEM[6143] = 8'h9B;
ROM_MEM[6144] = 8'hBA;
ROM_MEM[6145] = 8'h67;
ROM_MEM[6146] = 8'h62;
ROM_MEM[6147] = 8'h9B;
ROM_MEM[6148] = 8'h11;
ROM_MEM[6149] = 8'h80;
ROM_MEM[6150] = 8'hDA;
ROM_MEM[6151] = 8'h72;
ROM_MEM[6152] = 8'h04;
ROM_MEM[6153] = 8'h70;
ROM_MEM[6154] = 8'h99;
ROM_MEM[6155] = 8'hF5;
ROM_MEM[6156] = 8'h00;
ROM_MEM[6157] = 8'hCB;
ROM_MEM[6158] = 8'h09;
ROM_MEM[6159] = 8'hC0;
ROM_MEM[6160] = 8'h61;
ROM_MEM[6161] = 8'hC8;
ROM_MEM[6162] = 8'hCA;
ROM_MEM[6163] = 8'h42;
ROM_MEM[6164] = 8'h28;
ROM_MEM[6165] = 8'h9B;
ROM_MEM[6166] = 8'h94;
ROM_MEM[6167] = 8'hAE;
ROM_MEM[6168] = 8'h58;
ROM_MEM[6169] = 8'h69;
ROM_MEM[6170] = 8'hD0;
ROM_MEM[6171] = 8'h6A;
ROM_MEM[6172] = 8'hD2;
ROM_MEM[6173] = 8'hEA;
ROM_MEM[6174] = 8'h14;
ROM_MEM[6175] = 8'h35;
ROM_MEM[6176] = 8'h58;
ROM_MEM[6177] = 8'hCC;
ROM_MEM[6178] = 8'hED;
ROM_MEM[6179] = 8'hCA;
ROM_MEM[6180] = 8'h9B;
ROM_MEM[6181] = 8'h93;
ROM_MEM[6182] = 8'h21;
ROM_MEM[6183] = 8'hE1;
ROM_MEM[6184] = 8'hC5;
ROM_MEM[6185] = 8'h27;
ROM_MEM[6186] = 8'hCD;
ROM_MEM[6187] = 8'hDA;
ROM_MEM[6188] = 8'h5B;
ROM_MEM[6189] = 8'h84;
ROM_MEM[6190] = 8'h9E;
ROM_MEM[6191] = 8'h8E;
ROM_MEM[6192] = 8'h24;
ROM_MEM[6193] = 8'h19;
ROM_MEM[6194] = 8'h1F;
ROM_MEM[6195] = 8'h26;
ROM_MEM[6196] = 8'hBE;
ROM_MEM[6197] = 8'hDB;
ROM_MEM[6198] = 8'h32;
ROM_MEM[6199] = 8'hEF;
ROM_MEM[6200] = 8'h33;
ROM_MEM[6201] = 8'h49;
ROM_MEM[6202] = 8'h7C;
ROM_MEM[6203] = 8'h6E;
ROM_MEM[6204] = 8'hA8;
ROM_MEM[6205] = 8'h23;
ROM_MEM[6206] = 8'hCF;
ROM_MEM[6207] = 8'h54;
ROM_MEM[6208] = 8'hE5;
ROM_MEM[6209] = 8'hD8;
ROM_MEM[6210] = 8'hEE;
ROM_MEM[6211] = 8'h28;
ROM_MEM[6212] = 8'hDC;
ROM_MEM[6213] = 8'hD2;
ROM_MEM[6214] = 8'h48;
ROM_MEM[6215] = 8'h5C;
ROM_MEM[6216] = 8'h13;
ROM_MEM[6217] = 8'h80;
ROM_MEM[6218] = 8'h85;
ROM_MEM[6219] = 8'h2E;
ROM_MEM[6220] = 8'h04;
ROM_MEM[6221] = 8'h18;
ROM_MEM[6222] = 8'h9E;
ROM_MEM[6223] = 8'hA5;
ROM_MEM[6224] = 8'h80;
ROM_MEM[6225] = 8'hD4;
ROM_MEM[6226] = 8'h52;
ROM_MEM[6227] = 8'h15;
ROM_MEM[6228] = 8'h90;
ROM_MEM[6229] = 8'hB7;
ROM_MEM[6230] = 8'h0A;
ROM_MEM[6231] = 8'h01;
ROM_MEM[6232] = 8'h52;
ROM_MEM[6233] = 8'h15;
ROM_MEM[6234] = 8'h24;
ROM_MEM[6235] = 8'h40;
ROM_MEM[6236] = 8'hB4;
ROM_MEM[6237] = 8'h26;
ROM_MEM[6238] = 8'h04;
ROM_MEM[6239] = 8'h48;
ROM_MEM[6240] = 8'h5E;
ROM_MEM[6241] = 8'h19;
ROM_MEM[6242] = 8'h01;
ROM_MEM[6243] = 8'h9E;
ROM_MEM[6244] = 8'h85;
ROM_MEM[6245] = 8'h23;
ROM_MEM[6246] = 8'h40;
ROM_MEM[6247] = 8'h53;
ROM_MEM[6248] = 8'h73;
ROM_MEM[6249] = 8'h04;
ROM_MEM[6250] = 8'h78;
ROM_MEM[6251] = 8'h62;
ROM_MEM[6252] = 8'hC1;
ROM_MEM[6253] = 8'h80;
ROM_MEM[6254] = 8'hEA;
ROM_MEM[6255] = 8'h95;
ROM_MEM[6256] = 8'h0D;
ROM_MEM[6257] = 8'hD0;
ROM_MEM[6258] = 8'h82;
ROM_MEM[6259] = 8'h9B;
ROM_MEM[6260] = 8'h01;
ROM_MEM[6261] = 8'h6A;
ROM_MEM[6262] = 8'h74;
ROM_MEM[6263] = 8'h2B;
ROM_MEM[6264] = 8'h59;
ROM_MEM[6265] = 8'hA9;
ROM_MEM[6266] = 8'h1C;
ROM_MEM[6267] = 8'h2A;
ROM_MEM[6268] = 8'hDA;
ROM_MEM[6269] = 8'hE6;
ROM_MEM[6270] = 8'hA4;
ROM_MEM[6271] = 8'hB9;
ROM_MEM[6272] = 8'h68;
ROM_MEM[6273] = 8'h71;
ROM_MEM[6274] = 8'hEA;
ROM_MEM[6275] = 8'hA2;
ROM_MEM[6276] = 8'h93;
ROM_MEM[6277] = 8'hE4;
ROM_MEM[6278] = 8'h14;
ROM_MEM[6279] = 8'h45;
ROM_MEM[6280] = 8'hE9;
ROM_MEM[6281] = 8'hB5;
ROM_MEM[6282] = 8'h4F;
ROM_MEM[6283] = 8'h9C;
ROM_MEM[6284] = 8'h73;
ROM_MEM[6285] = 8'h04;
ROM_MEM[6286] = 8'hA7;
ROM_MEM[6287] = 8'h47;
ROM_MEM[6288] = 8'h5E;
ROM_MEM[6289] = 8'h49;
ROM_MEM[6290] = 8'h53;
ROM_MEM[6291] = 8'h61;
ROM_MEM[6292] = 8'hA6;
ROM_MEM[6293] = 8'h16;
ROM_MEM[6294] = 8'h79;
ROM_MEM[6295] = 8'hA7;
ROM_MEM[6296] = 8'h06;
ROM_MEM[6297] = 8'hB8;
ROM_MEM[6298] = 8'hD2;
ROM_MEM[6299] = 8'hDC;
ROM_MEM[6300] = 8'h00;
ROM_MEM[6301] = 8'h5B;
ROM_MEM[6302] = 8'h98;
ROM_MEM[6303] = 8'h2B;
ROM_MEM[6304] = 8'h60;
ROM_MEM[6305] = 8'h1B;
ROM_MEM[6306] = 8'h15;
ROM_MEM[6307] = 8'h50;
ROM_MEM[6308] = 8'h40;
ROM_MEM[6309] = 8'h73;
ROM_MEM[6310] = 8'h1A;
ROM_MEM[6311] = 8'hE0;
ROM_MEM[6312] = 8'hDA;
ROM_MEM[6313] = 8'hCA;
ROM_MEM[6314] = 8'hCD;
ROM_MEM[6315] = 8'hCC;
ROM_MEM[6316] = 8'hCC;
ROM_MEM[6317] = 8'h6E;
ROM_MEM[6318] = 8'hE9;
ROM_MEM[6319] = 8'hB3;
ROM_MEM[6320] = 8'h95;
ROM_MEM[6321] = 8'h30;
ROM_MEM[6322] = 8'hB5;
ROM_MEM[6323] = 8'hD8;
ROM_MEM[6324] = 8'hAB;
ROM_MEM[6325] = 8'hCF;
ROM_MEM[6326] = 8'h49;
ROM_MEM[6327] = 8'h5D;
ROM_MEM[6328] = 8'h22;
ROM_MEM[6329] = 8'h42;
ROM_MEM[6330] = 8'hAF;
ROM_MEM[6331] = 8'hA1;
ROM_MEM[6332] = 8'h56;
ROM_MEM[6333] = 8'h71;
ROM_MEM[6334] = 8'hAA;
ROM_MEM[6335] = 8'h34;
ROM_MEM[6336] = 8'hD3;
ROM_MEM[6337] = 8'h96;
ROM_MEM[6338] = 8'h9A;
ROM_MEM[6339] = 8'hC8;
ROM_MEM[6340] = 8'hAC;
ROM_MEM[6341] = 8'h42;
ROM_MEM[6342] = 8'h4A;
ROM_MEM[6343] = 8'hDB;
ROM_MEM[6344] = 8'h5A;
ROM_MEM[6345] = 8'h24;
ROM_MEM[6346] = 8'hE7;
ROM_MEM[6347] = 8'h4A;
ROM_MEM[6348] = 8'h39;
ROM_MEM[6349] = 8'h65;
ROM_MEM[6350] = 8'hEB;
ROM_MEM[6351] = 8'h8D;
ROM_MEM[6352] = 8'h42;
ROM_MEM[6353] = 8'h3B;
ROM_MEM[6354] = 8'hA4;
ROM_MEM[6355] = 8'hA4;
ROM_MEM[6356] = 8'hAD;
ROM_MEM[6357] = 8'h25;
ROM_MEM[6358] = 8'hB1;
ROM_MEM[6359] = 8'h48;
ROM_MEM[6360] = 8'h97;
ROM_MEM[6361] = 8'h8A;
ROM_MEM[6362] = 8'h80;
ROM_MEM[6363] = 8'h90;
ROM_MEM[6364] = 8'h62;
ROM_MEM[6365] = 8'h10;
ROM_MEM[6366] = 8'h10;
ROM_MEM[6367] = 8'h52;
ROM_MEM[6368] = 8'hF6;
ROM_MEM[6369] = 8'h03;
ROM_MEM[6370] = 8'h03;
ROM_MEM[6371] = 8'hB4;
ROM_MEM[6372] = 8'hE0;
ROM_MEM[6373] = 8'h59;
ROM_MEM[6374] = 8'h4B;
ROM_MEM[6375] = 8'h59;
ROM_MEM[6376] = 8'h4B;
ROM_MEM[6377] = 8'h59;
ROM_MEM[6378] = 8'h53;
ROM_MEM[6379] = 8'h59;
ROM_MEM[6380] = 8'h5B;
ROM_MEM[6381] = 8'h59;
ROM_MEM[6382] = 8'h63;
ROM_MEM[6383] = 8'h59;
ROM_MEM[6384] = 8'h6B;
ROM_MEM[6385] = 8'h59;
ROM_MEM[6386] = 8'h77;
ROM_MEM[6387] = 8'h59;
ROM_MEM[6388] = 8'h85;
ROM_MEM[6389] = 8'h59;
ROM_MEM[6390] = 8'hDD;
ROM_MEM[6391] = 8'h5A;
ROM_MEM[6392] = 8'h4B;
ROM_MEM[6393] = 8'h5A;
ROM_MEM[6394] = 8'hB9;
ROM_MEM[6395] = 8'h5D;
ROM_MEM[6396] = 8'h46;
ROM_MEM[6397] = 8'h5C;
ROM_MEM[6398] = 8'h7B;
ROM_MEM[6399] = 8'h5B;
ROM_MEM[6400] = 8'hCF;
ROM_MEM[6401] = 8'h5B;
ROM_MEM[6402] = 8'h27;
ROM_MEM[6403] = 8'h5E;
ROM_MEM[6404] = 8'h11;
ROM_MEM[6405] = 8'h5E;
ROM_MEM[6406] = 8'h97;
ROM_MEM[6407] = 8'h5F;
ROM_MEM[6408] = 8'h21;
ROM_MEM[6409] = 8'h5F;
ROM_MEM[6410] = 8'h95;
ROM_MEM[6411] = 8'h5F;
ROM_MEM[6412] = 8'hD5;
ROM_MEM[6413] = 8'h60;
ROM_MEM[6414] = 8'h37;
ROM_MEM[6415] = 8'h60;
ROM_MEM[6416] = 8'h99;
ROM_MEM[6417] = 8'h61;
ROM_MEM[6418] = 8'h49;
ROM_MEM[6419] = 8'h61;
ROM_MEM[6420] = 8'h8B;
ROM_MEM[6421] = 8'h62;
ROM_MEM[6422] = 8'h03;
ROM_MEM[6423] = 8'h62;
ROM_MEM[6424] = 8'h7B;
ROM_MEM[6425] = 8'h62;
ROM_MEM[6426] = 8'hF3;
ROM_MEM[6427] = 8'h63;
ROM_MEM[6428] = 8'h07;
ROM_MEM[6429] = 8'h63;
ROM_MEM[6430] = 8'h35;
ROM_MEM[6431] = 8'h63;
ROM_MEM[6432] = 8'h63;
ROM_MEM[6433] = 8'h63;
ROM_MEM[6434] = 8'h8D;
ROM_MEM[6435] = 8'h63;
ROM_MEM[6436] = 8'hB9;
ROM_MEM[6437] = 8'h64;
ROM_MEM[6438] = 8'h27;
ROM_MEM[6439] = 8'h64;
ROM_MEM[6440] = 8'hB1;
ROM_MEM[6441] = 8'h65;
ROM_MEM[6442] = 8'h4D;
ROM_MEM[6443] = 8'h65;
ROM_MEM[6444] = 8'hCB;
ROM_MEM[6445] = 8'h65;
ROM_MEM[6446] = 8'hFD;
ROM_MEM[6447] = 8'h66;
ROM_MEM[6448] = 8'h2B;
ROM_MEM[6449] = 8'h66;
ROM_MEM[6450] = 8'h3D;
ROM_MEM[6451] = 8'h66;
ROM_MEM[6452] = 8'h6B;
ROM_MEM[6453] = 8'h66;
ROM_MEM[6454] = 8'hB1;
ROM_MEM[6455] = 8'h66;
ROM_MEM[6456] = 8'hDD;
ROM_MEM[6457] = 8'h67;
ROM_MEM[6458] = 8'h07;
ROM_MEM[6459] = 8'h67;
ROM_MEM[6460] = 8'h43;
ROM_MEM[6461] = 8'h67;
ROM_MEM[6462] = 8'h75;
ROM_MEM[6463] = 8'h67;
ROM_MEM[6464] = 8'hA7;
ROM_MEM[6465] = 8'h67;
ROM_MEM[6466] = 8'hD3;
ROM_MEM[6467] = 8'h68;
ROM_MEM[6468] = 8'h07;
ROM_MEM[6469] = 8'h68;
ROM_MEM[6470] = 8'h0E;
ROM_MEM[6471] = 8'h68;
ROM_MEM[6472] = 8'h1D;
ROM_MEM[6473] = 8'h68;
ROM_MEM[6474] = 8'h2A;
ROM_MEM[6475] = 8'h8D;
ROM_MEM[6476] = 8'h06;
ROM_MEM[6477] = 8'h85;
ROM_MEM[6478] = 8'h00;
ROM_MEM[6479] = 8'h8D;
ROM_MEM[6480] = 8'h05;
ROM_MEM[6481] = 8'h00;
ROM_MEM[6482] = 8'h00;
ROM_MEM[6483] = 8'h8D;
ROM_MEM[6484] = 8'h06;
ROM_MEM[6485] = 8'h85;
ROM_MEM[6486] = 8'hFF;
ROM_MEM[6487] = 8'h8D;
ROM_MEM[6488] = 8'h05;
ROM_MEM[6489] = 8'h00;
ROM_MEM[6490] = 8'h00;
ROM_MEM[6491] = 8'h8D;
ROM_MEM[6492] = 8'h06;
ROM_MEM[6493] = 8'h85;
ROM_MEM[6494] = 8'hFD;
ROM_MEM[6495] = 8'h8D;
ROM_MEM[6496] = 8'h05;
ROM_MEM[6497] = 8'h00;
ROM_MEM[6498] = 8'h00;
ROM_MEM[6499] = 8'h8D;
ROM_MEM[6500] = 8'h06;
ROM_MEM[6501] = 8'h85;
ROM_MEM[6502] = 8'hFA;
ROM_MEM[6503] = 8'h8D;
ROM_MEM[6504] = 8'h05;
ROM_MEM[6505] = 8'h00;
ROM_MEM[6506] = 8'h00;
ROM_MEM[6507] = 8'h8E;
ROM_MEM[6508] = 8'h30;
ROM_MEM[6509] = 8'h41;
ROM_MEM[6510] = 8'h04;
ROM_MEM[6511] = 8'h85;
ROM_MEM[6512] = 8'hFF;
ROM_MEM[6513] = 8'h81;
ROM_MEM[6514] = 8'h01;
ROM_MEM[6515] = 8'h8F;
ROM_MEM[6516] = 8'h00;
ROM_MEM[6517] = 8'h00;
ROM_MEM[6518] = 8'h00;
ROM_MEM[6519] = 8'h84;
ROM_MEM[6520] = 8'h00;
ROM_MEM[6521] = 8'h82;
ROM_MEM[6522] = 8'h0F;
ROM_MEM[6523] = 8'h80;
ROM_MEM[6524] = 8'hCF;
ROM_MEM[6525] = 8'h8C;
ROM_MEM[6526] = 8'hFF;
ROM_MEM[6527] = 8'h8A;
ROM_MEM[6528] = 8'hA0;
ROM_MEM[6529] = 8'h87;
ROM_MEM[6530] = 8'h00;
ROM_MEM[6531] = 8'h00;
ROM_MEM[6532] = 8'h00;
ROM_MEM[6533] = 8'h80;
ROM_MEM[6534] = 8'h54;
ROM_MEM[6535] = 8'h87;
ROM_MEM[6536] = 8'h02;
ROM_MEM[6537] = 8'h33;
ROM_MEM[6538] = 8'h31;
ROM_MEM[6539] = 8'h33;
ROM_MEM[6540] = 8'h10;
ROM_MEM[6541] = 8'h38;
ROM_MEM[6542] = 8'h80;
ROM_MEM[6543] = 8'h3A;
ROM_MEM[6544] = 8'h40;
ROM_MEM[6545] = 8'h3A;
ROM_MEM[6546] = 8'h17;
ROM_MEM[6547] = 8'h3B;
ROM_MEM[6548] = 8'h16;
ROM_MEM[6549] = 8'h3D;
ROM_MEM[6550] = 8'h14;
ROM_MEM[6551] = 8'h3B;
ROM_MEM[6552] = 8'h80;
ROM_MEM[6553] = 8'h33;
ROM_MEM[6554] = 8'h40;
ROM_MEM[6555] = 8'h00;
ROM_MEM[6556] = 8'h20;
ROM_MEM[6557] = 8'h33;
ROM_MEM[6558] = 8'h20;
ROM_MEM[6559] = 8'h38;
ROM_MEM[6560] = 8'h60;
ROM_MEM[6561] = 8'h3A;
ROM_MEM[6562] = 8'h20;
ROM_MEM[6563] = 8'h3B;
ROM_MEM[6564] = 8'h20;
ROM_MEM[6565] = 8'h33;
ROM_MEM[6566] = 8'h20;
ROM_MEM[6567] = 8'h3B;
ROM_MEM[6568] = 8'h16;
ROM_MEM[6569] = 8'h38;
ROM_MEM[6570] = 8'h16;
ROM_MEM[6571] = 8'h3F;
ROM_MEM[6572] = 8'h14;
ROM_MEM[6573] = 8'h3D;
ROM_MEM[6574] = 8'hC0;
ROM_MEM[6575] = 8'h33;
ROM_MEM[6576] = 8'h30;
ROM_MEM[6577] = 8'h33;
ROM_MEM[6578] = 8'h10;
ROM_MEM[6579] = 8'h38;
ROM_MEM[6580] = 8'h40;
ROM_MEM[6581] = 8'h38;
ROM_MEM[6582] = 8'h31;
ROM_MEM[6583] = 8'h3A;
ROM_MEM[6584] = 8'h10;
ROM_MEM[6585] = 8'h3B;
ROM_MEM[6586] = 8'h30;
ROM_MEM[6587] = 8'h38;
ROM_MEM[6588] = 8'h10;
ROM_MEM[6589] = 8'h3F;
ROM_MEM[6590] = 8'h30;
ROM_MEM[6591] = 8'h3B;
ROM_MEM[6592] = 8'h10;
ROM_MEM[6593] = 8'h44;
ROM_MEM[6594] = 8'h80;
ROM_MEM[6595] = 8'h38;
ROM_MEM[6596] = 8'h40;
ROM_MEM[6597] = 8'h3B;
ROM_MEM[6598] = 8'h16;
ROM_MEM[6599] = 8'h3A;
ROM_MEM[6600] = 8'h16;
ROM_MEM[6601] = 8'h38;
ROM_MEM[6602] = 8'h14;
ROM_MEM[6603] = 8'h3F;
ROM_MEM[6604] = 8'h40;
ROM_MEM[6605] = 8'h3F;
ROM_MEM[6606] = 8'h17;
ROM_MEM[6607] = 8'h3B;
ROM_MEM[6608] = 8'h16;
ROM_MEM[6609] = 8'h38;
ROM_MEM[6610] = 8'h14;
ROM_MEM[6611] = 8'h33;
ROM_MEM[6612] = 8'h40;
ROM_MEM[6613] = 8'h33;
ROM_MEM[6614] = 8'h30;
ROM_MEM[6615] = 8'h33;
ROM_MEM[6616] = 8'h10;
ROM_MEM[6617] = 8'h38;
ROM_MEM[6618] = 8'hC0;
ROM_MEM[6619] = 8'h00;
ROM_MEM[6620] = 8'h00;
ROM_MEM[6621] = 8'h80;
ROM_MEM[6622] = 8'h54;
ROM_MEM[6623] = 8'h87;
ROM_MEM[6624] = 8'h03;
ROM_MEM[6625] = 8'h00;
ROM_MEM[6626] = 8'h40;
ROM_MEM[6627] = 8'h00;
ROM_MEM[6628] = 8'h40;
ROM_MEM[6629] = 8'h44;
ROM_MEM[6630] = 8'h20;
ROM_MEM[6631] = 8'h00;
ROM_MEM[6632] = 8'h40;
ROM_MEM[6633] = 8'h46;
ROM_MEM[6634] = 8'h20;
ROM_MEM[6635] = 8'h00;
ROM_MEM[6636] = 8'h20;
ROM_MEM[6637] = 8'h47;
ROM_MEM[6638] = 8'h20;
ROM_MEM[6639] = 8'h00;
ROM_MEM[6640] = 8'h40;
ROM_MEM[6641] = 8'h44;
ROM_MEM[6642] = 8'h20;
ROM_MEM[6643] = 8'h00;
ROM_MEM[6644] = 8'h40;
ROM_MEM[6645] = 8'h44;
ROM_MEM[6646] = 8'h20;
ROM_MEM[6647] = 8'h43;
ROM_MEM[6648] = 8'h16;
ROM_MEM[6649] = 8'h43;
ROM_MEM[6650] = 8'h16;
ROM_MEM[6651] = 8'h43;
ROM_MEM[6652] = 8'h14;
ROM_MEM[6653] = 8'h00;
ROM_MEM[6654] = 8'h40;
ROM_MEM[6655] = 8'h44;
ROM_MEM[6656] = 8'h20;
ROM_MEM[6657] = 8'h00;
ROM_MEM[6658] = 8'h40;
ROM_MEM[6659] = 8'h47;
ROM_MEM[6660] = 8'h20;
ROM_MEM[6661] = 8'h00;
ROM_MEM[6662] = 8'h20;
ROM_MEM[6663] = 8'h47;
ROM_MEM[6664] = 8'h20;
ROM_MEM[6665] = 8'h00;
ROM_MEM[6666] = 8'h40;
ROM_MEM[6667] = 8'h44;
ROM_MEM[6668] = 8'h16;
ROM_MEM[6669] = 8'h44;
ROM_MEM[6670] = 8'h16;
ROM_MEM[6671] = 8'h44;
ROM_MEM[6672] = 8'h14;
ROM_MEM[6673] = 8'h44;
ROM_MEM[6674] = 8'h21;
ROM_MEM[6675] = 8'h44;
ROM_MEM[6676] = 8'h20;
ROM_MEM[6677] = 8'h46;
ROM_MEM[6678] = 8'h20;
ROM_MEM[6679] = 8'h46;
ROM_MEM[6680] = 8'h20;
ROM_MEM[6681] = 8'h00;
ROM_MEM[6682] = 8'h40;
ROM_MEM[6683] = 8'h44;
ROM_MEM[6684] = 8'h20;
ROM_MEM[6685] = 8'h00;
ROM_MEM[6686] = 8'h40;
ROM_MEM[6687] = 8'h44;
ROM_MEM[6688] = 8'h20;
ROM_MEM[6689] = 8'h00;
ROM_MEM[6690] = 8'h20;
ROM_MEM[6691] = 8'h44;
ROM_MEM[6692] = 8'h20;
ROM_MEM[6693] = 8'h00;
ROM_MEM[6694] = 8'h40;
ROM_MEM[6695] = 8'h47;
ROM_MEM[6696] = 8'h20;
ROM_MEM[6697] = 8'h47;
ROM_MEM[6698] = 8'h20;
ROM_MEM[6699] = 8'h47;
ROM_MEM[6700] = 8'h20;
ROM_MEM[6701] = 8'h47;
ROM_MEM[6702] = 8'h20;
ROM_MEM[6703] = 8'h47;
ROM_MEM[6704] = 8'h16;
ROM_MEM[6705] = 8'h47;
ROM_MEM[6706] = 8'h16;
ROM_MEM[6707] = 8'h47;
ROM_MEM[6708] = 8'h14;
ROM_MEM[6709] = 8'h00;
ROM_MEM[6710] = 8'h40;
ROM_MEM[6711] = 8'h47;
ROM_MEM[6712] = 8'h20;
ROM_MEM[6713] = 8'h00;
ROM_MEM[6714] = 8'h40;
ROM_MEM[6715] = 8'h46;
ROM_MEM[6716] = 8'h20;
ROM_MEM[6717] = 8'h00;
ROM_MEM[6718] = 8'h20;
ROM_MEM[6719] = 8'h46;
ROM_MEM[6720] = 8'h20;
ROM_MEM[6721] = 8'h00;
ROM_MEM[6722] = 8'h40;
ROM_MEM[6723] = 8'h44;
ROM_MEM[6724] = 8'h20;
ROM_MEM[6725] = 8'h44;
ROM_MEM[6726] = 8'h20;
ROM_MEM[6727] = 8'h44;
ROM_MEM[6728] = 8'h40;
ROM_MEM[6729] = 8'h00;
ROM_MEM[6730] = 8'h00;
ROM_MEM[6731] = 8'h80;
ROM_MEM[6732] = 8'h54;
ROM_MEM[6733] = 8'h87;
ROM_MEM[6734] = 8'h03;
ROM_MEM[6735] = 8'h00;
ROM_MEM[6736] = 8'h40;
ROM_MEM[6737] = 8'h00;
ROM_MEM[6738] = 8'h40;
ROM_MEM[6739] = 8'h3B;
ROM_MEM[6740] = 8'h20;
ROM_MEM[6741] = 8'h00;
ROM_MEM[6742] = 8'h40;
ROM_MEM[6743] = 8'h3F;
ROM_MEM[6744] = 8'h20;
ROM_MEM[6745] = 8'h00;
ROM_MEM[6746] = 8'h20;
ROM_MEM[6747] = 8'h43;
ROM_MEM[6748] = 8'h20;
ROM_MEM[6749] = 8'h00;
ROM_MEM[6750] = 8'h40;
ROM_MEM[6751] = 8'h3F;
ROM_MEM[6752] = 8'h20;
ROM_MEM[6753] = 8'h00;
ROM_MEM[6754] = 8'h40;
ROM_MEM[6755] = 8'h3B;
ROM_MEM[6756] = 8'h20;
ROM_MEM[6757] = 8'h3A;
ROM_MEM[6758] = 8'h16;
ROM_MEM[6759] = 8'h3A;
ROM_MEM[6760] = 8'h16;
ROM_MEM[6761] = 8'h3A;
ROM_MEM[6762] = 8'h14;
ROM_MEM[6763] = 8'h00;
ROM_MEM[6764] = 8'h40;
ROM_MEM[6765] = 8'h3B;
ROM_MEM[6766] = 8'h20;
ROM_MEM[6767] = 8'h00;
ROM_MEM[6768] = 8'h40;
ROM_MEM[6769] = 8'h3F;
ROM_MEM[6770] = 8'h20;
ROM_MEM[6771] = 8'h00;
ROM_MEM[6772] = 8'h20;
ROM_MEM[6773] = 8'h3F;
ROM_MEM[6774] = 8'h20;
ROM_MEM[6775] = 8'h00;
ROM_MEM[6776] = 8'h40;
ROM_MEM[6777] = 8'h41;
ROM_MEM[6778] = 8'h16;
ROM_MEM[6779] = 8'h41;
ROM_MEM[6780] = 8'h16;
ROM_MEM[6781] = 8'h41;
ROM_MEM[6782] = 8'h14;
ROM_MEM[6783] = 8'h41;
ROM_MEM[6784] = 8'h21;
ROM_MEM[6785] = 8'h41;
ROM_MEM[6786] = 8'h20;
ROM_MEM[6787] = 8'h43;
ROM_MEM[6788] = 8'h20;
ROM_MEM[6789] = 8'h43;
ROM_MEM[6790] = 8'h20;
ROM_MEM[6791] = 8'h00;
ROM_MEM[6792] = 8'h40;
ROM_MEM[6793] = 8'h3B;
ROM_MEM[6794] = 8'h20;
ROM_MEM[6795] = 8'h00;
ROM_MEM[6796] = 8'h40;
ROM_MEM[6797] = 8'h3F;
ROM_MEM[6798] = 8'h20;
ROM_MEM[6799] = 8'h00;
ROM_MEM[6800] = 8'h20;
ROM_MEM[6801] = 8'h3B;
ROM_MEM[6802] = 8'h20;
ROM_MEM[6803] = 8'h00;
ROM_MEM[6804] = 8'h40;
ROM_MEM[6805] = 8'h40;
ROM_MEM[6806] = 8'h20;
ROM_MEM[6807] = 8'h40;
ROM_MEM[6808] = 8'h20;
ROM_MEM[6809] = 8'h40;
ROM_MEM[6810] = 8'h20;
ROM_MEM[6811] = 8'h40;
ROM_MEM[6812] = 8'h20;
ROM_MEM[6813] = 8'h40;
ROM_MEM[6814] = 8'h16;
ROM_MEM[6815] = 8'h40;
ROM_MEM[6816] = 8'h16;
ROM_MEM[6817] = 8'h40;
ROM_MEM[6818] = 8'h14;
ROM_MEM[6819] = 8'h00;
ROM_MEM[6820] = 8'h40;
ROM_MEM[6821] = 8'h44;
ROM_MEM[6822] = 8'h20;
ROM_MEM[6823] = 8'h00;
ROM_MEM[6824] = 8'h40;
ROM_MEM[6825] = 8'h44;
ROM_MEM[6826] = 8'h20;
ROM_MEM[6827] = 8'h00;
ROM_MEM[6828] = 8'h20;
ROM_MEM[6829] = 8'h43;
ROM_MEM[6830] = 8'h20;
ROM_MEM[6831] = 8'h00;
ROM_MEM[6832] = 8'h40;
ROM_MEM[6833] = 8'h3B;
ROM_MEM[6834] = 8'h20;
ROM_MEM[6835] = 8'h3B;
ROM_MEM[6836] = 8'h20;
ROM_MEM[6837] = 8'h3B;
ROM_MEM[6838] = 8'h40;
ROM_MEM[6839] = 8'h00;
ROM_MEM[6840] = 8'h00;
ROM_MEM[6841] = 8'h80;
ROM_MEM[6842] = 8'h54;
ROM_MEM[6843] = 8'h87;
ROM_MEM[6844] = 8'h03;
ROM_MEM[6845] = 8'h00;
ROM_MEM[6846] = 8'h40;
ROM_MEM[6847] = 8'h00;
ROM_MEM[6848] = 8'h40;
ROM_MEM[6849] = 8'h20;
ROM_MEM[6850] = 8'h20;
ROM_MEM[6851] = 8'h00;
ROM_MEM[6852] = 8'h40;
ROM_MEM[6853] = 8'h20;
ROM_MEM[6854] = 8'h20;
ROM_MEM[6855] = 8'h00;
ROM_MEM[6856] = 8'h20;
ROM_MEM[6857] = 8'h20;
ROM_MEM[6858] = 8'h20;
ROM_MEM[6859] = 8'h00;
ROM_MEM[6860] = 8'h40;
ROM_MEM[6861] = 8'h20;
ROM_MEM[6862] = 8'h20;
ROM_MEM[6863] = 8'h00;
ROM_MEM[6864] = 8'h40;
ROM_MEM[6865] = 8'h20;
ROM_MEM[6866] = 8'h20;
ROM_MEM[6867] = 8'h1B;
ROM_MEM[6868] = 8'h16;
ROM_MEM[6869] = 8'h1B;
ROM_MEM[6870] = 8'h16;
ROM_MEM[6871] = 8'h1B;
ROM_MEM[6872] = 8'h14;
ROM_MEM[6873] = 8'h00;
ROM_MEM[6874] = 8'h40;
ROM_MEM[6875] = 8'h20;
ROM_MEM[6876] = 8'h20;
ROM_MEM[6877] = 8'h00;
ROM_MEM[6878] = 8'h40;
ROM_MEM[6879] = 8'h20;
ROM_MEM[6880] = 8'h20;
ROM_MEM[6881] = 8'h00;
ROM_MEM[6882] = 8'h20;
ROM_MEM[6883] = 8'h20;
ROM_MEM[6884] = 8'h20;
ROM_MEM[6885] = 8'h00;
ROM_MEM[6886] = 8'h40;
ROM_MEM[6887] = 8'h19;
ROM_MEM[6888] = 8'h16;
ROM_MEM[6889] = 8'h19;
ROM_MEM[6890] = 8'h16;
ROM_MEM[6891] = 8'h19;
ROM_MEM[6892] = 8'h14;
ROM_MEM[6893] = 8'h19;
ROM_MEM[6894] = 8'h21;
ROM_MEM[6895] = 8'h19;
ROM_MEM[6896] = 8'h20;
ROM_MEM[6897] = 8'h1B;
ROM_MEM[6898] = 8'h20;
ROM_MEM[6899] = 8'h1B;
ROM_MEM[6900] = 8'h20;
ROM_MEM[6901] = 8'h00;
ROM_MEM[6902] = 8'h40;
ROM_MEM[6903] = 8'h20;
ROM_MEM[6904] = 8'h20;
ROM_MEM[6905] = 8'h00;
ROM_MEM[6906] = 8'h40;
ROM_MEM[6907] = 8'h20;
ROM_MEM[6908] = 8'h20;
ROM_MEM[6909] = 8'h00;
ROM_MEM[6910] = 8'h20;
ROM_MEM[6911] = 8'h20;
ROM_MEM[6912] = 8'h20;
ROM_MEM[6913] = 8'h00;
ROM_MEM[6914] = 8'h40;
ROM_MEM[6915] = 8'h1C;
ROM_MEM[6916] = 8'h20;
ROM_MEM[6917] = 8'h1C;
ROM_MEM[6918] = 8'h20;
ROM_MEM[6919] = 8'h1C;
ROM_MEM[6920] = 8'h20;
ROM_MEM[6921] = 8'h1C;
ROM_MEM[6922] = 8'h20;
ROM_MEM[6923] = 8'h1C;
ROM_MEM[6924] = 8'h16;
ROM_MEM[6925] = 8'h1C;
ROM_MEM[6926] = 8'h16;
ROM_MEM[6927] = 8'h1C;
ROM_MEM[6928] = 8'h14;
ROM_MEM[6929] = 8'h00;
ROM_MEM[6930] = 8'h40;
ROM_MEM[6931] = 8'h1B;
ROM_MEM[6932] = 8'h20;
ROM_MEM[6933] = 8'h00;
ROM_MEM[6934] = 8'h40;
ROM_MEM[6935] = 8'h1B;
ROM_MEM[6936] = 8'h20;
ROM_MEM[6937] = 8'h00;
ROM_MEM[6938] = 8'h20;
ROM_MEM[6939] = 8'h1B;
ROM_MEM[6940] = 8'h20;
ROM_MEM[6941] = 8'h00;
ROM_MEM[6942] = 8'h40;
ROM_MEM[6943] = 8'h20;
ROM_MEM[6944] = 8'h20;
ROM_MEM[6945] = 8'h20;
ROM_MEM[6946] = 8'h20;
ROM_MEM[6947] = 8'h20;
ROM_MEM[6948] = 8'h40;
ROM_MEM[6949] = 8'h00;
ROM_MEM[6950] = 8'h00;
ROM_MEM[6951] = 8'h80;
ROM_MEM[6952] = 8'h96;
ROM_MEM[6953] = 8'h87;
ROM_MEM[6954] = 8'h01;
ROM_MEM[6955] = 8'h82;
ROM_MEM[6956] = 8'h07;
ROM_MEM[6957] = 8'h8E;
ROM_MEM[6958] = 8'h02;
ROM_MEM[6959] = 8'h90;
ROM_MEM[6960] = 8'h5B;
ROM_MEM[6961] = 8'hAC;
ROM_MEM[6962] = 8'h8F;
ROM_MEM[6963] = 8'h00;
ROM_MEM[6964] = 8'h27;
ROM_MEM[6965] = 8'h40;
ROM_MEM[6966] = 8'h00;
ROM_MEM[6967] = 8'h40;
ROM_MEM[6968] = 8'h25;
ROM_MEM[6969] = 8'h40;
ROM_MEM[6970] = 8'h00;
ROM_MEM[6971] = 8'h40;
ROM_MEM[6972] = 8'h90;
ROM_MEM[6973] = 8'h5B;
ROM_MEM[6974] = 8'hB5;
ROM_MEM[6975] = 8'h8E;
ROM_MEM[6976] = 8'h02;
ROM_MEM[6977] = 8'h90;
ROM_MEM[6978] = 8'h5B;
ROM_MEM[6979] = 8'hAC;
ROM_MEM[6980] = 8'h8F;
ROM_MEM[6981] = 8'h00;
ROM_MEM[6982] = 8'h20;
ROM_MEM[6983] = 8'h40;
ROM_MEM[6984] = 8'h00;
ROM_MEM[6985] = 8'h40;
ROM_MEM[6986] = 8'h20;
ROM_MEM[6987] = 8'h40;
ROM_MEM[6988] = 8'h00;
ROM_MEM[6989] = 8'h40;
ROM_MEM[6990] = 8'h25;
ROM_MEM[6991] = 8'h40;
ROM_MEM[6992] = 8'h27;
ROM_MEM[6993] = 8'h40;
ROM_MEM[6994] = 8'h28;
ROM_MEM[6995] = 8'h40;
ROM_MEM[6996] = 8'h29;
ROM_MEM[6997] = 8'h40;
ROM_MEM[6998] = 8'h8E;
ROM_MEM[6999] = 8'h02;
ROM_MEM[7000] = 8'h90;
ROM_MEM[7001] = 8'h5B;
ROM_MEM[7002] = 8'hAC;
ROM_MEM[7003] = 8'h8F;
ROM_MEM[7004] = 8'h00;
ROM_MEM[7005] = 8'h25;
ROM_MEM[7006] = 8'h40;
ROM_MEM[7007] = 8'h00;
ROM_MEM[7008] = 8'h40;
ROM_MEM[7009] = 8'h25;
ROM_MEM[7010] = 8'h40;
ROM_MEM[7011] = 8'h00;
ROM_MEM[7012] = 8'h40;
ROM_MEM[7013] = 8'h90;
ROM_MEM[7014] = 8'h5B;
ROM_MEM[7015] = 8'hB5;
ROM_MEM[7016] = 8'h23;
ROM_MEM[7017] = 8'h40;
ROM_MEM[7018] = 8'h00;
ROM_MEM[7019] = 8'h40;
ROM_MEM[7020] = 8'h23;
ROM_MEM[7021] = 8'h40;
ROM_MEM[7022] = 8'h00;
ROM_MEM[7023] = 8'h40;
ROM_MEM[7024] = 8'h2A;
ROM_MEM[7025] = 8'h40;
ROM_MEM[7026] = 8'h00;
ROM_MEM[7027] = 8'h40;
ROM_MEM[7028] = 8'h27;
ROM_MEM[7029] = 8'h40;
ROM_MEM[7030] = 8'h00;
ROM_MEM[7031] = 8'h40;
ROM_MEM[7032] = 8'h2C;
ROM_MEM[7033] = 8'h40;
ROM_MEM[7034] = 8'h00;
ROM_MEM[7035] = 8'h40;
ROM_MEM[7036] = 8'h25;
ROM_MEM[7037] = 8'h40;
ROM_MEM[7038] = 8'h00;
ROM_MEM[7039] = 8'h40;
ROM_MEM[7040] = 8'h2A;
ROM_MEM[7041] = 8'h40;
ROM_MEM[7042] = 8'h29;
ROM_MEM[7043] = 8'h40;
ROM_MEM[7044] = 8'h27;
ROM_MEM[7045] = 8'h40;
ROM_MEM[7046] = 8'h25;
ROM_MEM[7047] = 8'h40;
ROM_MEM[7048] = 8'h8E;
ROM_MEM[7049] = 8'h03;
ROM_MEM[7050] = 8'h90;
ROM_MEM[7051] = 8'h5B;
ROM_MEM[7052] = 8'hBE;
ROM_MEM[7053] = 8'h8F;
ROM_MEM[7054] = 8'h00;
ROM_MEM[7055] = 8'h27;
ROM_MEM[7056] = 8'h20;
ROM_MEM[7057] = 8'h00;
ROM_MEM[7058] = 8'h20;
ROM_MEM[7059] = 8'h00;
ROM_MEM[7060] = 8'hC0;
ROM_MEM[7061] = 8'h00;
ROM_MEM[7062] = 8'hC0;
ROM_MEM[7063] = 8'h22;
ROM_MEM[7064] = 8'h40;
ROM_MEM[7065] = 8'h8E;
ROM_MEM[7066] = 8'h03;
ROM_MEM[7067] = 8'h90;
ROM_MEM[7068] = 8'h5B;
ROM_MEM[7069] = 8'hBE;
ROM_MEM[7070] = 8'h8F;
ROM_MEM[7071] = 8'h00;
ROM_MEM[7072] = 8'h27;
ROM_MEM[7073] = 8'h40;
ROM_MEM[7074] = 8'h23;
ROM_MEM[7075] = 8'h40;
ROM_MEM[7076] = 8'h22;
ROM_MEM[7077] = 8'h40;
ROM_MEM[7078] = 8'h22;
ROM_MEM[7079] = 8'h20;
ROM_MEM[7080] = 8'h27;
ROM_MEM[7081] = 8'h40;
ROM_MEM[7082] = 8'h00;
ROM_MEM[7083] = 8'h00;
ROM_MEM[7084] = 8'h27;
ROM_MEM[7085] = 8'h40;
ROM_MEM[7086] = 8'h00;
ROM_MEM[7087] = 8'h40;
ROM_MEM[7088] = 8'h22;
ROM_MEM[7089] = 8'h40;
ROM_MEM[7090] = 8'h00;
ROM_MEM[7091] = 8'h40;
ROM_MEM[7092] = 8'h91;
ROM_MEM[7093] = 8'h2A;
ROM_MEM[7094] = 8'h40;
ROM_MEM[7095] = 8'h00;
ROM_MEM[7096] = 8'h40;
ROM_MEM[7097] = 8'h25;
ROM_MEM[7098] = 8'h40;
ROM_MEM[7099] = 8'h00;
ROM_MEM[7100] = 8'h40;
ROM_MEM[7101] = 8'h91;
ROM_MEM[7102] = 8'h27;
ROM_MEM[7103] = 8'h40;
ROM_MEM[7104] = 8'h25;
ROM_MEM[7105] = 8'h40;
ROM_MEM[7106] = 8'h23;
ROM_MEM[7107] = 8'h40;
ROM_MEM[7108] = 8'h22;
ROM_MEM[7109] = 8'h40;
ROM_MEM[7110] = 8'h20;
ROM_MEM[7111] = 8'h40;
ROM_MEM[7112] = 8'h1E;
ROM_MEM[7113] = 8'h40;
ROM_MEM[7114] = 8'h1D;
ROM_MEM[7115] = 8'h40;
ROM_MEM[7116] = 8'h1B;
ROM_MEM[7117] = 8'h40;
ROM_MEM[7118] = 8'h91;
ROM_MEM[7119] = 8'h80;
ROM_MEM[7120] = 8'h96;
ROM_MEM[7121] = 8'h87;
ROM_MEM[7122] = 8'h01;
ROM_MEM[7123] = 8'h82;
ROM_MEM[7124] = 8'h03;
ROM_MEM[7125] = 8'h90;
ROM_MEM[7126] = 8'h5C;
ROM_MEM[7127] = 8'h6A;
ROM_MEM[7128] = 8'h33;
ROM_MEM[7129] = 8'h20;
ROM_MEM[7130] = 8'h33;
ROM_MEM[7131] = 8'h40;
ROM_MEM[7132] = 8'h33;
ROM_MEM[7133] = 8'h20;
ROM_MEM[7134] = 8'h32;
ROM_MEM[7135] = 8'h20;
ROM_MEM[7136] = 8'h33;
ROM_MEM[7137] = 8'h20;
ROM_MEM[7138] = 8'h31;
ROM_MEM[7139] = 8'h20;
ROM_MEM[7140] = 8'h00;
ROM_MEM[7141] = 8'h20;
ROM_MEM[7142] = 8'h30;
ROM_MEM[7143] = 8'h20;
ROM_MEM[7144] = 8'h31;
ROM_MEM[7145] = 8'h20;
ROM_MEM[7146] = 8'h2F;
ROM_MEM[7147] = 8'h20;
ROM_MEM[7148] = 8'h2E;
ROM_MEM[7149] = 8'h60;
ROM_MEM[7150] = 8'h2A;
ROM_MEM[7151] = 8'h20;
ROM_MEM[7152] = 8'h2A;
ROM_MEM[7153] = 8'h81;
ROM_MEM[7154] = 8'h90;
ROM_MEM[7155] = 8'h5C;
ROM_MEM[7156] = 8'h6A;
ROM_MEM[7157] = 8'h32;
ROM_MEM[7158] = 8'h20;
ROM_MEM[7159] = 8'h33;
ROM_MEM[7160] = 8'h40;
ROM_MEM[7161] = 8'h30;
ROM_MEM[7162] = 8'h20;
ROM_MEM[7163] = 8'h00;
ROM_MEM[7164] = 8'h20;
ROM_MEM[7165] = 8'h30;
ROM_MEM[7166] = 8'h40;
ROM_MEM[7167] = 8'h30;
ROM_MEM[7168] = 8'h21;
ROM_MEM[7169] = 8'h2F;
ROM_MEM[7170] = 8'h20;
ROM_MEM[7171] = 8'h30;
ROM_MEM[7172] = 8'h40;
ROM_MEM[7173] = 8'h35;
ROM_MEM[7174] = 8'h20;
ROM_MEM[7175] = 8'h33;
ROM_MEM[7176] = 8'h40;
ROM_MEM[7177] = 8'h31;
ROM_MEM[7178] = 8'h40;
ROM_MEM[7179] = 8'h2F;
ROM_MEM[7180] = 8'h60;
ROM_MEM[7181] = 8'h90;
ROM_MEM[7182] = 8'h5C;
ROM_MEM[7183] = 8'h6A;
ROM_MEM[7184] = 8'h33;
ROM_MEM[7185] = 8'h20;
ROM_MEM[7186] = 8'h33;
ROM_MEM[7187] = 8'h40;
ROM_MEM[7188] = 8'h35;
ROM_MEM[7189] = 8'h20;
ROM_MEM[7190] = 8'h00;
ROM_MEM[7191] = 8'h20;
ROM_MEM[7192] = 8'h35;
ROM_MEM[7193] = 8'h40;
ROM_MEM[7194] = 8'h35;
ROM_MEM[7195] = 8'h21;
ROM_MEM[7196] = 8'h31;
ROM_MEM[7197] = 8'h20;
ROM_MEM[7198] = 8'h2F;
ROM_MEM[7199] = 8'h40;
ROM_MEM[7200] = 8'h2D;
ROM_MEM[7201] = 8'h60;
ROM_MEM[7202] = 8'h2A;
ROM_MEM[7203] = 8'h20;
ROM_MEM[7204] = 8'h2A;
ROM_MEM[7205] = 8'h81;
ROM_MEM[7206] = 8'h8C;
ROM_MEM[7207] = 8'hFF;
ROM_MEM[7208] = 8'h87;
ROM_MEM[7209] = 8'h04;
ROM_MEM[7210] = 8'h2A;
ROM_MEM[7211] = 8'h80;
ROM_MEM[7212] = 8'h2F;
ROM_MEM[7213] = 8'h81;
ROM_MEM[7214] = 8'h31;
ROM_MEM[7215] = 8'h81;
ROM_MEM[7216] = 8'h37;
ROM_MEM[7217] = 8'h81;
ROM_MEM[7218] = 8'h8C;
ROM_MEM[7219] = 8'h00;
ROM_MEM[7220] = 8'h87;
ROM_MEM[7221] = 8'h01;
ROM_MEM[7222] = 8'h38;
ROM_MEM[7223] = 8'h40;
ROM_MEM[7224] = 8'h37;
ROM_MEM[7225] = 8'h40;
ROM_MEM[7226] = 8'h30;
ROM_MEM[7227] = 8'h20;
ROM_MEM[7228] = 8'h2F;
ROM_MEM[7229] = 8'h40;
ROM_MEM[7230] = 8'h2E;
ROM_MEM[7231] = 8'h20;
ROM_MEM[7232] = 8'h00;
ROM_MEM[7233] = 8'h80;
ROM_MEM[7234] = 8'h00;
ROM_MEM[7235] = 8'h81;
ROM_MEM[7236] = 8'h8E;
ROM_MEM[7237] = 8'h10;
ROM_MEM[7238] = 8'h00;
ROM_MEM[7239] = 8'h80;
ROM_MEM[7240] = 8'h8F;
ROM_MEM[7241] = 8'h00;
ROM_MEM[7242] = 8'h8E;
ROM_MEM[7243] = 8'h03;
ROM_MEM[7244] = 8'h00;
ROM_MEM[7245] = 8'h40;
ROM_MEM[7246] = 8'h33;
ROM_MEM[7247] = 8'hC0;
ROM_MEM[7248] = 8'h33;
ROM_MEM[7249] = 8'h81;
ROM_MEM[7250] = 8'h32;
ROM_MEM[7251] = 8'h20;
ROM_MEM[7252] = 8'h00;
ROM_MEM[7253] = 8'h60;
ROM_MEM[7254] = 8'h8F;
ROM_MEM[7255] = 8'h00;
ROM_MEM[7256] = 8'h86;
ROM_MEM[7257] = 8'h01;
ROM_MEM[7258] = 8'h00;
ROM_MEM[7259] = 8'h20;
ROM_MEM[7260] = 8'h33;
ROM_MEM[7261] = 8'h20;
ROM_MEM[7262] = 8'h00;
ROM_MEM[7263] = 8'h20;
ROM_MEM[7264] = 8'h33;
ROM_MEM[7265] = 8'h20;
ROM_MEM[7266] = 8'h00;
ROM_MEM[7267] = 8'h60;
ROM_MEM[7268] = 8'h33;
ROM_MEM[7269] = 8'h40;
ROM_MEM[7270] = 8'h86;
ROM_MEM[7271] = 8'h00;
ROM_MEM[7272] = 8'h00;
ROM_MEM[7273] = 8'h00;
ROM_MEM[7274] = 8'h33;
ROM_MEM[7275] = 8'h40;
ROM_MEM[7276] = 8'h36;
ROM_MEM[7277] = 8'h40;
ROM_MEM[7278] = 8'h33;
ROM_MEM[7279] = 8'h40;
ROM_MEM[7280] = 8'h36;
ROM_MEM[7281] = 8'h40;
ROM_MEM[7282] = 8'h33;
ROM_MEM[7283] = 8'h20;
ROM_MEM[7284] = 8'h36;
ROM_MEM[7285] = 8'h41;
ROM_MEM[7286] = 8'h33;
ROM_MEM[7287] = 8'h20;
ROM_MEM[7288] = 8'h00;
ROM_MEM[7289] = 8'h20;
ROM_MEM[7290] = 8'h91;
ROM_MEM[7291] = 8'h80;
ROM_MEM[7292] = 8'h96;
ROM_MEM[7293] = 8'h87;
ROM_MEM[7294] = 8'h01;
ROM_MEM[7295] = 8'h82;
ROM_MEM[7296] = 8'h03;
ROM_MEM[7297] = 8'h90;
ROM_MEM[7298] = 8'h5D;
ROM_MEM[7299] = 8'h16;
ROM_MEM[7300] = 8'h36;
ROM_MEM[7301] = 8'h20;
ROM_MEM[7302] = 8'h35;
ROM_MEM[7303] = 8'h20;
ROM_MEM[7304] = 8'h36;
ROM_MEM[7305] = 8'h20;
ROM_MEM[7306] = 8'h35;
ROM_MEM[7307] = 8'h20;
ROM_MEM[7308] = 8'h00;
ROM_MEM[7309] = 8'h20;
ROM_MEM[7310] = 8'h34;
ROM_MEM[7311] = 8'h20;
ROM_MEM[7312] = 8'h35;
ROM_MEM[7313] = 8'h20;
ROM_MEM[7314] = 8'h32;
ROM_MEM[7315] = 8'h20;
ROM_MEM[7316] = 8'h31;
ROM_MEM[7317] = 8'h60;
ROM_MEM[7318] = 8'h2E;
ROM_MEM[7319] = 8'h20;
ROM_MEM[7320] = 8'h2E;
ROM_MEM[7321] = 8'h81;
ROM_MEM[7322] = 8'h90;
ROM_MEM[7323] = 8'h5D;
ROM_MEM[7324] = 8'h16;
ROM_MEM[7325] = 8'h33;
ROM_MEM[7326] = 8'h20;
ROM_MEM[7327] = 8'h00;
ROM_MEM[7328] = 8'h20;
ROM_MEM[7329] = 8'h33;
ROM_MEM[7330] = 8'h40;
ROM_MEM[7331] = 8'h33;
ROM_MEM[7332] = 8'h21;
ROM_MEM[7333] = 8'h32;
ROM_MEM[7334] = 8'h20;
ROM_MEM[7335] = 8'h33;
ROM_MEM[7336] = 8'h40;
ROM_MEM[7337] = 8'h38;
ROM_MEM[7338] = 8'h20;
ROM_MEM[7339] = 8'h36;
ROM_MEM[7340] = 8'h40;
ROM_MEM[7341] = 8'h35;
ROM_MEM[7342] = 8'h40;
ROM_MEM[7343] = 8'h33;
ROM_MEM[7344] = 8'h60;
ROM_MEM[7345] = 8'h90;
ROM_MEM[7346] = 8'h5D;
ROM_MEM[7347] = 8'h16;
ROM_MEM[7348] = 8'h38;
ROM_MEM[7349] = 8'h20;
ROM_MEM[7350] = 8'h00;
ROM_MEM[7351] = 8'h20;
ROM_MEM[7352] = 8'h38;
ROM_MEM[7353] = 8'h40;
ROM_MEM[7354] = 8'h38;
ROM_MEM[7355] = 8'h21;
ROM_MEM[7356] = 8'h35;
ROM_MEM[7357] = 8'h20;
ROM_MEM[7358] = 8'h35;
ROM_MEM[7359] = 8'h40;
ROM_MEM[7360] = 8'h31;
ROM_MEM[7361] = 8'h60;
ROM_MEM[7362] = 8'h2E;
ROM_MEM[7363] = 8'h20;
ROM_MEM[7364] = 8'h2E;
ROM_MEM[7365] = 8'h81;
ROM_MEM[7366] = 8'h8C;
ROM_MEM[7367] = 8'hFF;
ROM_MEM[7368] = 8'h87;
ROM_MEM[7369] = 8'h04;
ROM_MEM[7370] = 8'h2F;
ROM_MEM[7371] = 8'h80;
ROM_MEM[7372] = 8'h33;
ROM_MEM[7373] = 8'h81;
ROM_MEM[7374] = 8'h36;
ROM_MEM[7375] = 8'h81;
ROM_MEM[7376] = 8'h3A;
ROM_MEM[7377] = 8'h81;
ROM_MEM[7378] = 8'h8C;
ROM_MEM[7379] = 8'h00;
ROM_MEM[7380] = 8'h87;
ROM_MEM[7381] = 8'h01;
ROM_MEM[7382] = 8'h3B;
ROM_MEM[7383] = 8'h40;
ROM_MEM[7384] = 8'h3A;
ROM_MEM[7385] = 8'h40;
ROM_MEM[7386] = 8'h35;
ROM_MEM[7387] = 8'h20;
ROM_MEM[7388] = 8'h31;
ROM_MEM[7389] = 8'h41;
ROM_MEM[7390] = 8'h31;
ROM_MEM[7391] = 8'h20;
ROM_MEM[7392] = 8'h00;
ROM_MEM[7393] = 8'h80;
ROM_MEM[7394] = 8'h00;
ROM_MEM[7395] = 8'h81;
ROM_MEM[7396] = 8'h8E;
ROM_MEM[7397] = 8'h03;
ROM_MEM[7398] = 8'h90;
ROM_MEM[7399] = 8'h5D;
ROM_MEM[7400] = 8'h2B;
ROM_MEM[7401] = 8'h8F;
ROM_MEM[7402] = 8'h00;
ROM_MEM[7403] = 8'h00;
ROM_MEM[7404] = 8'h20;
ROM_MEM[7405] = 8'h8E;
ROM_MEM[7406] = 8'h03;
ROM_MEM[7407] = 8'h33;
ROM_MEM[7408] = 8'h20;
ROM_MEM[7409] = 8'h36;
ROM_MEM[7410] = 8'h20;
ROM_MEM[7411] = 8'h33;
ROM_MEM[7412] = 8'h20;
ROM_MEM[7413] = 8'h35;
ROM_MEM[7414] = 8'h20;
ROM_MEM[7415] = 8'h8F;
ROM_MEM[7416] = 8'h00;
ROM_MEM[7417] = 8'h33;
ROM_MEM[7418] = 8'h20;
ROM_MEM[7419] = 8'h36;
ROM_MEM[7420] = 8'h20;
ROM_MEM[7421] = 8'h00;
ROM_MEM[7422] = 8'h20;
ROM_MEM[7423] = 8'h8E;
ROM_MEM[7424] = 8'h03;
ROM_MEM[7425] = 8'h90;
ROM_MEM[7426] = 8'h5D;
ROM_MEM[7427] = 8'h2B;
ROM_MEM[7428] = 8'h8F;
ROM_MEM[7429] = 8'h00;
ROM_MEM[7430] = 8'h33;
ROM_MEM[7431] = 8'h20;
ROM_MEM[7432] = 8'h33;
ROM_MEM[7433] = 8'h20;
ROM_MEM[7434] = 8'h36;
ROM_MEM[7435] = 8'h20;
ROM_MEM[7436] = 8'h33;
ROM_MEM[7437] = 8'h20;
ROM_MEM[7438] = 8'h36;
ROM_MEM[7439] = 8'h20;
ROM_MEM[7440] = 8'h36;
ROM_MEM[7441] = 8'h40;
ROM_MEM[7442] = 8'h33;
ROM_MEM[7443] = 8'h40;
ROM_MEM[7444] = 8'h00;
ROM_MEM[7445] = 8'h00;
ROM_MEM[7446] = 8'h36;
ROM_MEM[7447] = 8'h40;
ROM_MEM[7448] = 8'h3A;
ROM_MEM[7449] = 8'h40;
ROM_MEM[7450] = 8'h36;
ROM_MEM[7451] = 8'h40;
ROM_MEM[7452] = 8'h3A;
ROM_MEM[7453] = 8'h40;
ROM_MEM[7454] = 8'h36;
ROM_MEM[7455] = 8'h20;
ROM_MEM[7456] = 8'h3A;
ROM_MEM[7457] = 8'h41;
ROM_MEM[7458] = 8'h36;
ROM_MEM[7459] = 8'h20;
ROM_MEM[7460] = 8'h00;
ROM_MEM[7461] = 8'h20;
ROM_MEM[7462] = 8'h35;
ROM_MEM[7463] = 8'h20;
ROM_MEM[7464] = 8'h36;
ROM_MEM[7465] = 8'h40;
ROM_MEM[7466] = 8'h91;
ROM_MEM[7467] = 8'h33;
ROM_MEM[7468] = 8'h40;
ROM_MEM[7469] = 8'h00;
ROM_MEM[7470] = 8'h20;
ROM_MEM[7471] = 8'h36;
ROM_MEM[7472] = 8'h40;
ROM_MEM[7473] = 8'h33;
ROM_MEM[7474] = 8'h20;
ROM_MEM[7475] = 8'h35;
ROM_MEM[7476] = 8'h40;
ROM_MEM[7477] = 8'h00;
ROM_MEM[7478] = 8'h20;
ROM_MEM[7479] = 8'h33;
ROM_MEM[7480] = 8'h20;
ROM_MEM[7481] = 8'h36;
ROM_MEM[7482] = 8'h20;
ROM_MEM[7483] = 8'h33;
ROM_MEM[7484] = 8'h20;
ROM_MEM[7485] = 8'h35;
ROM_MEM[7486] = 8'h20;
ROM_MEM[7487] = 8'h33;
ROM_MEM[7488] = 8'h20;
ROM_MEM[7489] = 8'h36;
ROM_MEM[7490] = 8'h20;
ROM_MEM[7491] = 8'h00;
ROM_MEM[7492] = 8'h20;
ROM_MEM[7493] = 8'h91;
ROM_MEM[7494] = 8'h80;
ROM_MEM[7495] = 8'h96;
ROM_MEM[7496] = 8'h87;
ROM_MEM[7497] = 8'h01;
ROM_MEM[7498] = 8'h82;
ROM_MEM[7499] = 8'h03;
ROM_MEM[7500] = 8'h90;
ROM_MEM[7501] = 8'h5D;
ROM_MEM[7502] = 8'hE1;
ROM_MEM[7503] = 8'h3A;
ROM_MEM[7504] = 8'h20;
ROM_MEM[7505] = 8'h39;
ROM_MEM[7506] = 8'h20;
ROM_MEM[7507] = 8'h3A;
ROM_MEM[7508] = 8'h20;
ROM_MEM[7509] = 8'h38;
ROM_MEM[7510] = 8'h20;
ROM_MEM[7511] = 8'h00;
ROM_MEM[7512] = 8'h20;
ROM_MEM[7513] = 8'h37;
ROM_MEM[7514] = 8'h20;
ROM_MEM[7515] = 8'h38;
ROM_MEM[7516] = 8'h20;
ROM_MEM[7517] = 8'h37;
ROM_MEM[7518] = 8'h20;
ROM_MEM[7519] = 8'h36;
ROM_MEM[7520] = 8'h60;
ROM_MEM[7521] = 8'h33;
ROM_MEM[7522] = 8'h20;
ROM_MEM[7523] = 8'h33;
ROM_MEM[7524] = 8'h81;
ROM_MEM[7525] = 8'h90;
ROM_MEM[7526] = 8'h5D;
ROM_MEM[7527] = 8'hE1;
ROM_MEM[7528] = 8'h38;
ROM_MEM[7529] = 8'h20;
ROM_MEM[7530] = 8'h00;
ROM_MEM[7531] = 8'h20;
ROM_MEM[7532] = 8'h38;
ROM_MEM[7533] = 8'h40;
ROM_MEM[7534] = 8'h38;
ROM_MEM[7535] = 8'h21;
ROM_MEM[7536] = 8'h37;
ROM_MEM[7537] = 8'h20;
ROM_MEM[7538] = 8'h38;
ROM_MEM[7539] = 8'h40;
ROM_MEM[7540] = 8'h3D;
ROM_MEM[7541] = 8'h20;
ROM_MEM[7542] = 8'h3B;
ROM_MEM[7543] = 8'h40;
ROM_MEM[7544] = 8'h3A;
ROM_MEM[7545] = 8'h40;
ROM_MEM[7546] = 8'h38;
ROM_MEM[7547] = 8'h60;
ROM_MEM[7548] = 8'h90;
ROM_MEM[7549] = 8'h5D;
ROM_MEM[7550] = 8'hE1;
ROM_MEM[7551] = 8'h3D;
ROM_MEM[7552] = 8'h20;
ROM_MEM[7553] = 8'h00;
ROM_MEM[7554] = 8'h20;
ROM_MEM[7555] = 8'h3D;
ROM_MEM[7556] = 8'h40;
ROM_MEM[7557] = 8'h3D;
ROM_MEM[7558] = 8'h21;
ROM_MEM[7559] = 8'h3A;
ROM_MEM[7560] = 8'h20;
ROM_MEM[7561] = 8'h38;
ROM_MEM[7562] = 8'h40;
ROM_MEM[7563] = 8'h36;
ROM_MEM[7564] = 8'h60;
ROM_MEM[7565] = 8'h33;
ROM_MEM[7566] = 8'h20;
ROM_MEM[7567] = 8'h33;
ROM_MEM[7568] = 8'h81;
ROM_MEM[7569] = 8'h8C;
ROM_MEM[7570] = 8'hFF;
ROM_MEM[7571] = 8'h87;
ROM_MEM[7572] = 8'h04;
ROM_MEM[7573] = 8'h33;
ROM_MEM[7574] = 8'h80;
ROM_MEM[7575] = 8'h36;
ROM_MEM[7576] = 8'h81;
ROM_MEM[7577] = 8'h3A;
ROM_MEM[7578] = 8'h81;
ROM_MEM[7579] = 8'h3D;
ROM_MEM[7580] = 8'h81;
ROM_MEM[7581] = 8'h8C;
ROM_MEM[7582] = 8'h00;
ROM_MEM[7583] = 8'h87;
ROM_MEM[7584] = 8'h01;
ROM_MEM[7585] = 8'h40;
ROM_MEM[7586] = 8'h41;
ROM_MEM[7587] = 8'h3F;
ROM_MEM[7588] = 8'h40;
ROM_MEM[7589] = 8'h39;
ROM_MEM[7590] = 8'h20;
ROM_MEM[7591] = 8'h3A;
ROM_MEM[7592] = 8'h41;
ROM_MEM[7593] = 8'h36;
ROM_MEM[7594] = 8'h20;
ROM_MEM[7595] = 8'h00;
ROM_MEM[7596] = 8'h80;
ROM_MEM[7597] = 8'h00;
ROM_MEM[7598] = 8'h81;
ROM_MEM[7599] = 8'h8E;
ROM_MEM[7600] = 8'h03;
ROM_MEM[7601] = 8'h90;
ROM_MEM[7602] = 8'h5D;
ROM_MEM[7603] = 8'hF6;
ROM_MEM[7604] = 8'h8F;
ROM_MEM[7605] = 8'h00;
ROM_MEM[7606] = 8'h36;
ROM_MEM[7607] = 8'h20;
ROM_MEM[7608] = 8'h8E;
ROM_MEM[7609] = 8'h03;
ROM_MEM[7610] = 8'h36;
ROM_MEM[7611] = 8'h20;
ROM_MEM[7612] = 8'h39;
ROM_MEM[7613] = 8'h20;
ROM_MEM[7614] = 8'h36;
ROM_MEM[7615] = 8'h20;
ROM_MEM[7616] = 8'h38;
ROM_MEM[7617] = 8'h20;
ROM_MEM[7618] = 8'h8F;
ROM_MEM[7619] = 8'h00;
ROM_MEM[7620] = 8'h36;
ROM_MEM[7621] = 8'h20;
ROM_MEM[7622] = 8'h39;
ROM_MEM[7623] = 8'h20;
ROM_MEM[7624] = 8'h33;
ROM_MEM[7625] = 8'h20;
ROM_MEM[7626] = 8'h8E;
ROM_MEM[7627] = 8'h03;
ROM_MEM[7628] = 8'h90;
ROM_MEM[7629] = 8'h5D;
ROM_MEM[7630] = 8'hF6;
ROM_MEM[7631] = 8'h8F;
ROM_MEM[7632] = 8'h00;
ROM_MEM[7633] = 8'h36;
ROM_MEM[7634] = 8'h20;
ROM_MEM[7635] = 8'h36;
ROM_MEM[7636] = 8'h20;
ROM_MEM[7637] = 8'h39;
ROM_MEM[7638] = 8'h20;
ROM_MEM[7639] = 8'h36;
ROM_MEM[7640] = 8'h20;
ROM_MEM[7641] = 8'h39;
ROM_MEM[7642] = 8'h20;
ROM_MEM[7643] = 8'h39;
ROM_MEM[7644] = 8'h40;
ROM_MEM[7645] = 8'h36;
ROM_MEM[7646] = 8'h40;
ROM_MEM[7647] = 8'h00;
ROM_MEM[7648] = 8'h00;
ROM_MEM[7649] = 8'h3A;
ROM_MEM[7650] = 8'h40;
ROM_MEM[7651] = 8'h3F;
ROM_MEM[7652] = 8'h40;
ROM_MEM[7653] = 8'h3A;
ROM_MEM[7654] = 8'h40;
ROM_MEM[7655] = 8'h3F;
ROM_MEM[7656] = 8'h40;
ROM_MEM[7657] = 8'h3A;
ROM_MEM[7658] = 8'h20;
ROM_MEM[7659] = 8'h3F;
ROM_MEM[7660] = 8'h41;
ROM_MEM[7661] = 8'h3A;
ROM_MEM[7662] = 8'h20;
ROM_MEM[7663] = 8'h00;
ROM_MEM[7664] = 8'h20;
ROM_MEM[7665] = 8'h39;
ROM_MEM[7666] = 8'h20;
ROM_MEM[7667] = 8'h3A;
ROM_MEM[7668] = 8'h40;
ROM_MEM[7669] = 8'h91;
ROM_MEM[7670] = 8'h36;
ROM_MEM[7671] = 8'h40;
ROM_MEM[7672] = 8'h00;
ROM_MEM[7673] = 8'h20;
ROM_MEM[7674] = 8'h39;
ROM_MEM[7675] = 8'h40;
ROM_MEM[7676] = 8'h36;
ROM_MEM[7677] = 8'h20;
ROM_MEM[7678] = 8'h38;
ROM_MEM[7679] = 8'h40;
ROM_MEM[7680] = 8'h00;
ROM_MEM[7681] = 8'h20;
ROM_MEM[7682] = 8'h36;
ROM_MEM[7683] = 8'h20;
ROM_MEM[7684] = 8'h39;
ROM_MEM[7685] = 8'h20;
ROM_MEM[7686] = 8'h36;
ROM_MEM[7687] = 8'h20;
ROM_MEM[7688] = 8'h38;
ROM_MEM[7689] = 8'h20;
ROM_MEM[7690] = 8'h36;
ROM_MEM[7691] = 8'h20;
ROM_MEM[7692] = 8'h39;
ROM_MEM[7693] = 8'h20;
ROM_MEM[7694] = 8'h33;
ROM_MEM[7695] = 8'h20;
ROM_MEM[7696] = 8'h91;
ROM_MEM[7697] = 8'h80;
ROM_MEM[7698] = 8'h80;
ROM_MEM[7699] = 8'h87;
ROM_MEM[7700] = 8'h02;
ROM_MEM[7701] = 8'h84;
ROM_MEM[7702] = 8'h0C;
ROM_MEM[7703] = 8'h82;
ROM_MEM[7704] = 8'h05;
ROM_MEM[7705] = 8'h00;
ROM_MEM[7706] = 8'h80;
ROM_MEM[7707] = 8'h4F;
ROM_MEM[7708] = 8'h20;
ROM_MEM[7709] = 8'h47;
ROM_MEM[7710] = 8'h20;
ROM_MEM[7711] = 8'h4E;
ROM_MEM[7712] = 8'h20;
ROM_MEM[7713] = 8'h4D;
ROM_MEM[7714] = 8'h20;
ROM_MEM[7715] = 8'h4A;
ROM_MEM[7716] = 8'h20;
ROM_MEM[7717] = 8'h42;
ROM_MEM[7718] = 8'h20;
ROM_MEM[7719] = 8'h49;
ROM_MEM[7720] = 8'h20;
ROM_MEM[7721] = 8'h47;
ROM_MEM[7722] = 8'h20;
ROM_MEM[7723] = 8'h46;
ROM_MEM[7724] = 8'h20;
ROM_MEM[7725] = 8'h3D;
ROM_MEM[7726] = 8'h20;
ROM_MEM[7727] = 8'h43;
ROM_MEM[7728] = 8'h20;
ROM_MEM[7729] = 8'h42;
ROM_MEM[7730] = 8'h20;
ROM_MEM[7731] = 8'h3D;
ROM_MEM[7732] = 8'h20;
ROM_MEM[7733] = 8'h36;
ROM_MEM[7734] = 8'h20;
ROM_MEM[7735] = 8'h3E;
ROM_MEM[7736] = 8'h20;
ROM_MEM[7737] = 8'h3D;
ROM_MEM[7738] = 8'h20;
ROM_MEM[7739] = 8'h8E;
ROM_MEM[7740] = 8'h02;
ROM_MEM[7741] = 8'h43;
ROM_MEM[7742] = 8'h20;
ROM_MEM[7743] = 8'h3B;
ROM_MEM[7744] = 8'h20;
ROM_MEM[7745] = 8'h42;
ROM_MEM[7746] = 8'h20;
ROM_MEM[7747] = 8'h41;
ROM_MEM[7748] = 8'h20;
ROM_MEM[7749] = 8'h3E;
ROM_MEM[7750] = 8'h20;
ROM_MEM[7751] = 8'h36;
ROM_MEM[7752] = 8'h20;
ROM_MEM[7753] = 8'h3B;
ROM_MEM[7754] = 8'h20;
ROM_MEM[7755] = 8'h3A;
ROM_MEM[7756] = 8'h20;
ROM_MEM[7757] = 8'h8F;
ROM_MEM[7758] = 8'h00;
ROM_MEM[7759] = 8'h84;
ROM_MEM[7760] = 8'h00;
ROM_MEM[7761] = 8'h82;
ROM_MEM[7762] = 8'h0A;
ROM_MEM[7763] = 8'h3E;
ROM_MEM[7764] = 8'h80;
ROM_MEM[7765] = 8'h42;
ROM_MEM[7766] = 8'h80;
ROM_MEM[7767] = 8'h82;
ROM_MEM[7768] = 8'h09;
ROM_MEM[7769] = 8'h87;
ROM_MEM[7770] = 8'h03;
ROM_MEM[7771] = 8'h8E;
ROM_MEM[7772] = 8'h04;
ROM_MEM[7773] = 8'h3E;
ROM_MEM[7774] = 8'h40;
ROM_MEM[7775] = 8'h8F;
ROM_MEM[7776] = 8'h00;
ROM_MEM[7777] = 8'h48;
ROM_MEM[7778] = 8'h80;
ROM_MEM[7779] = 8'h48;
ROM_MEM[7780] = 8'h81;
ROM_MEM[7781] = 8'h47;
ROM_MEM[7782] = 8'hC0;
ROM_MEM[7783] = 8'h47;
ROM_MEM[7784] = 8'h40;
ROM_MEM[7785] = 8'h45;
ROM_MEM[7786] = 8'h60;
ROM_MEM[7787] = 8'h45;
ROM_MEM[7788] = 8'h11;
ROM_MEM[7789] = 8'h82;
ROM_MEM[7790] = 8'h07;
ROM_MEM[7791] = 8'h44;
ROM_MEM[7792] = 8'h0C;
ROM_MEM[7793] = 8'h00;
ROM_MEM[7794] = 8'h04;
ROM_MEM[7795] = 8'h8E;
ROM_MEM[7796] = 8'h03;
ROM_MEM[7797] = 8'h44;
ROM_MEM[7798] = 8'h40;
ROM_MEM[7799] = 8'h41;
ROM_MEM[7800] = 8'h10;
ROM_MEM[7801] = 8'h00;
ROM_MEM[7802] = 8'h20;
ROM_MEM[7803] = 8'h44;
ROM_MEM[7804] = 8'h0C;
ROM_MEM[7805] = 8'h00;
ROM_MEM[7806] = 8'h04;
ROM_MEM[7807] = 8'h8F;
ROM_MEM[7808] = 8'h00;
ROM_MEM[7809] = 8'h87;
ROM_MEM[7810] = 8'h02;
ROM_MEM[7811] = 8'h45;
ROM_MEM[7812] = 8'hC0;
ROM_MEM[7813] = 8'h45;
ROM_MEM[7814] = 8'hC1;
ROM_MEM[7815] = 8'h45;
ROM_MEM[7816] = 8'h81;
ROM_MEM[7817] = 8'h83;
ROM_MEM[7818] = 8'hFF;
ROM_MEM[7819] = 8'h45;
ROM_MEM[7820] = 8'h41;
ROM_MEM[7821] = 8'h83;
ROM_MEM[7822] = 8'hFF;
ROM_MEM[7823] = 8'h45;
ROM_MEM[7824] = 8'h41;
ROM_MEM[7825] = 8'h83;
ROM_MEM[7826] = 8'hFF;
ROM_MEM[7827] = 8'h45;
ROM_MEM[7828] = 8'h41;
ROM_MEM[7829] = 8'h00;
ROM_MEM[7830] = 8'h00;
ROM_MEM[7831] = 8'h80;
ROM_MEM[7832] = 8'h80;
ROM_MEM[7833] = 8'h87;
ROM_MEM[7834] = 8'h03;
ROM_MEM[7835] = 8'h84;
ROM_MEM[7836] = 8'h0C;
ROM_MEM[7837] = 8'h82;
ROM_MEM[7838] = 8'h05;
ROM_MEM[7839] = 8'h00;
ROM_MEM[7840] = 8'h80;
ROM_MEM[7841] = 8'h43;
ROM_MEM[7842] = 8'h40;
ROM_MEM[7843] = 8'h42;
ROM_MEM[7844] = 8'h20;
ROM_MEM[7845] = 8'h41;
ROM_MEM[7846] = 8'h20;
ROM_MEM[7847] = 8'h3E;
ROM_MEM[7848] = 8'h40;
ROM_MEM[7849] = 8'h3D;
ROM_MEM[7850] = 8'h20;
ROM_MEM[7851] = 8'h3B;
ROM_MEM[7852] = 8'h20;
ROM_MEM[7853] = 8'h3A;
ROM_MEM[7854] = 8'h40;
ROM_MEM[7855] = 8'h37;
ROM_MEM[7856] = 8'h20;
ROM_MEM[7857] = 8'h36;
ROM_MEM[7858] = 8'h20;
ROM_MEM[7859] = 8'h31;
ROM_MEM[7860] = 8'h40;
ROM_MEM[7861] = 8'h32;
ROM_MEM[7862] = 8'h20;
ROM_MEM[7863] = 8'h31;
ROM_MEM[7864] = 8'h20;
ROM_MEM[7865] = 8'h37;
ROM_MEM[7866] = 8'h40;
ROM_MEM[7867] = 8'h36;
ROM_MEM[7868] = 8'h20;
ROM_MEM[7869] = 8'h35;
ROM_MEM[7870] = 8'h20;
ROM_MEM[7871] = 8'h32;
ROM_MEM[7872] = 8'h40;
ROM_MEM[7873] = 8'h3B;
ROM_MEM[7874] = 8'h20;
ROM_MEM[7875] = 8'h3A;
ROM_MEM[7876] = 8'h20;
ROM_MEM[7877] = 8'h37;
ROM_MEM[7878] = 8'h40;
ROM_MEM[7879] = 8'h36;
ROM_MEM[7880] = 8'h40;
ROM_MEM[7881] = 8'h32;
ROM_MEM[7882] = 8'h40;
ROM_MEM[7883] = 8'h00;
ROM_MEM[7884] = 8'h40;
ROM_MEM[7885] = 8'h84;
ROM_MEM[7886] = 8'h00;
ROM_MEM[7887] = 8'h87;
ROM_MEM[7888] = 8'h02;
ROM_MEM[7889] = 8'h82;
ROM_MEM[7890] = 8'h0A;
ROM_MEM[7891] = 8'h3B;
ROM_MEM[7892] = 8'h80;
ROM_MEM[7893] = 8'h32;
ROM_MEM[7894] = 8'h20;
ROM_MEM[7895] = 8'h36;
ROM_MEM[7896] = 8'h20;
ROM_MEM[7897] = 8'h3B;
ROM_MEM[7898] = 8'h16;
ROM_MEM[7899] = 8'h3E;
ROM_MEM[7900] = 8'h16;
ROM_MEM[7901] = 8'h42;
ROM_MEM[7902] = 8'h14;
ROM_MEM[7903] = 8'h82;
ROM_MEM[7904] = 8'h09;
ROM_MEM[7905] = 8'h87;
ROM_MEM[7906] = 8'h03;
ROM_MEM[7907] = 8'h8E;
ROM_MEM[7908] = 8'h04;
ROM_MEM[7909] = 8'h45;
ROM_MEM[7910] = 8'h40;
ROM_MEM[7911] = 8'h8F;
ROM_MEM[7912] = 8'h00;
ROM_MEM[7913] = 8'h45;
ROM_MEM[7914] = 8'h80;
ROM_MEM[7915] = 8'h45;
ROM_MEM[7916] = 8'h81;
ROM_MEM[7917] = 8'h44;
ROM_MEM[7918] = 8'hC0;
ROM_MEM[7919] = 8'h44;
ROM_MEM[7920] = 8'h40;
ROM_MEM[7921] = 8'h42;
ROM_MEM[7922] = 8'h80;
ROM_MEM[7923] = 8'h42;
ROM_MEM[7924] = 8'h81;
ROM_MEM[7925] = 8'h42;
ROM_MEM[7926] = 8'h81;
ROM_MEM[7927] = 8'h42;
ROM_MEM[7928] = 8'h81;
ROM_MEM[7929] = 8'h82;
ROM_MEM[7930] = 8'h07;
ROM_MEM[7931] = 8'h00;
ROM_MEM[7932] = 8'h80;
ROM_MEM[7933] = 8'h1A;
ROM_MEM[7934] = 8'h40;
ROM_MEM[7935] = 8'h21;
ROM_MEM[7936] = 8'h40;
ROM_MEM[7937] = 8'h2A;
ROM_MEM[7938] = 8'h40;
ROM_MEM[7939] = 8'h2D;
ROM_MEM[7940] = 8'h40;
ROM_MEM[7941] = 8'h32;
ROM_MEM[7942] = 8'h20;
ROM_MEM[7943] = 8'h39;
ROM_MEM[7944] = 8'h20;
ROM_MEM[7945] = 8'h3E;
ROM_MEM[7946] = 8'h16;
ROM_MEM[7947] = 8'h86;
ROM_MEM[7948] = 8'h01;
ROM_MEM[7949] = 8'h42;
ROM_MEM[7950] = 8'h16;
ROM_MEM[7951] = 8'h45;
ROM_MEM[7952] = 8'h14;
ROM_MEM[7953] = 8'h86;
ROM_MEM[7954] = 8'h00;
ROM_MEM[7955] = 8'h83;
ROM_MEM[7956] = 8'hFF;
ROM_MEM[7957] = 8'h4A;
ROM_MEM[7958] = 8'h40;
ROM_MEM[7959] = 8'h83;
ROM_MEM[7960] = 8'hFF;
ROM_MEM[7961] = 8'h4A;
ROM_MEM[7962] = 8'h41;
ROM_MEM[7963] = 8'h83;
ROM_MEM[7964] = 8'hFF;
ROM_MEM[7965] = 8'h4A;
ROM_MEM[7966] = 8'h41;
ROM_MEM[7967] = 8'h00;
ROM_MEM[7968] = 8'h00;
ROM_MEM[7969] = 8'h80;
ROM_MEM[7970] = 8'h80;
ROM_MEM[7971] = 8'h87;
ROM_MEM[7972] = 8'h03;
ROM_MEM[7973] = 8'h82;
ROM_MEM[7974] = 8'h05;
ROM_MEM[7975] = 8'h00;
ROM_MEM[7976] = 8'h10;
ROM_MEM[7977] = 8'h86;
ROM_MEM[7978] = 8'h01;
ROM_MEM[7979] = 8'h25;
ROM_MEM[7980] = 8'h10;
ROM_MEM[7981] = 8'h86;
ROM_MEM[7982] = 8'h00;
ROM_MEM[7983] = 8'h26;
ROM_MEM[7984] = 8'h10;
ROM_MEM[7985] = 8'h29;
ROM_MEM[7986] = 8'h10;
ROM_MEM[7987] = 8'h2A;
ROM_MEM[7988] = 8'h10;
ROM_MEM[7989] = 8'h2C;
ROM_MEM[7990] = 8'h10;
ROM_MEM[7991] = 8'h2E;
ROM_MEM[7992] = 8'h10;
ROM_MEM[7993] = 8'h2F;
ROM_MEM[7994] = 8'h10;
ROM_MEM[7995] = 8'h4F;
ROM_MEM[7996] = 8'h40;
ROM_MEM[7997] = 8'h00;
ROM_MEM[7998] = 8'hC0;
ROM_MEM[7999] = 8'h8E;
ROM_MEM[8000] = 8'h06;
ROM_MEM[8001] = 8'h00;
ROM_MEM[8002] = 8'h80;
ROM_MEM[8003] = 8'h8F;
ROM_MEM[8004] = 8'h00;
ROM_MEM[8005] = 8'h87;
ROM_MEM[8006] = 8'h02;
ROM_MEM[8007] = 8'h82;
ROM_MEM[8008] = 8'h0A;
ROM_MEM[8009] = 8'h36;
ROM_MEM[8010] = 8'h80;
ROM_MEM[8011] = 8'h2F;
ROM_MEM[8012] = 8'h20;
ROM_MEM[8013] = 8'h32;
ROM_MEM[8014] = 8'h20;
ROM_MEM[8015] = 8'h36;
ROM_MEM[8016] = 8'h16;
ROM_MEM[8017] = 8'h3B;
ROM_MEM[8018] = 8'h16;
ROM_MEM[8019] = 8'h3E;
ROM_MEM[8020] = 8'h14;
ROM_MEM[8021] = 8'h82;
ROM_MEM[8022] = 8'h09;
ROM_MEM[8023] = 8'h87;
ROM_MEM[8024] = 8'h03;
ROM_MEM[8025] = 8'h8E;
ROM_MEM[8026] = 8'h04;
ROM_MEM[8027] = 8'h42;
ROM_MEM[8028] = 8'h40;
ROM_MEM[8029] = 8'h8F;
ROM_MEM[8030] = 8'h00;
ROM_MEM[8031] = 8'h41;
ROM_MEM[8032] = 8'h80;
ROM_MEM[8033] = 8'h41;
ROM_MEM[8034] = 8'h81;
ROM_MEM[8035] = 8'h40;
ROM_MEM[8036] = 8'hC0;
ROM_MEM[8037] = 8'h40;
ROM_MEM[8038] = 8'h40;
ROM_MEM[8039] = 8'h00;
ROM_MEM[8040] = 8'h40;
ROM_MEM[8041] = 8'h00;
ROM_MEM[8042] = 8'h30;
ROM_MEM[8043] = 8'h82;
ROM_MEM[8044] = 8'h07;
ROM_MEM[8045] = 8'h41;
ROM_MEM[8046] = 8'h0C;
ROM_MEM[8047] = 8'h00;
ROM_MEM[8048] = 8'h04;
ROM_MEM[8049] = 8'h8E;
ROM_MEM[8050] = 8'h03;
ROM_MEM[8051] = 8'h41;
ROM_MEM[8052] = 8'h40;
ROM_MEM[8053] = 8'h3E;
ROM_MEM[8054] = 8'h10;
ROM_MEM[8055] = 8'h00;
ROM_MEM[8056] = 8'h20;
ROM_MEM[8057] = 8'h41;
ROM_MEM[8058] = 8'h0C;
ROM_MEM[8059] = 8'h00;
ROM_MEM[8060] = 8'h04;
ROM_MEM[8061] = 8'h8F;
ROM_MEM[8062] = 8'h00;
ROM_MEM[8063] = 8'h87;
ROM_MEM[8064] = 8'h02;
ROM_MEM[8065] = 8'h42;
ROM_MEM[8066] = 8'hC0;
ROM_MEM[8067] = 8'h42;
ROM_MEM[8068] = 8'hC1;
ROM_MEM[8069] = 8'h42;
ROM_MEM[8070] = 8'h81;
ROM_MEM[8071] = 8'h83;
ROM_MEM[8072] = 8'hFF;
ROM_MEM[8073] = 8'h42;
ROM_MEM[8074] = 8'h41;
ROM_MEM[8075] = 8'h83;
ROM_MEM[8076] = 8'hFF;
ROM_MEM[8077] = 8'h42;
ROM_MEM[8078] = 8'h41;
ROM_MEM[8079] = 8'h83;
ROM_MEM[8080] = 8'hFF;
ROM_MEM[8081] = 8'h42;
ROM_MEM[8082] = 8'h41;
ROM_MEM[8083] = 8'h00;
ROM_MEM[8084] = 8'h00;
ROM_MEM[8085] = 8'h80;
ROM_MEM[8086] = 8'h80;
ROM_MEM[8087] = 8'h87;
ROM_MEM[8088] = 8'h02;
ROM_MEM[8089] = 8'h82;
ROM_MEM[8090] = 8'h05;
ROM_MEM[8091] = 8'h25;
ROM_MEM[8092] = 8'hC0;
ROM_MEM[8093] = 8'h25;
ROM_MEM[8094] = 8'hC1;
ROM_MEM[8095] = 8'h25;
ROM_MEM[8096] = 8'hC1;
ROM_MEM[8097] = 8'h25;
ROM_MEM[8098] = 8'hC1;
ROM_MEM[8099] = 8'h25;
ROM_MEM[8100] = 8'hC1;
ROM_MEM[8101] = 8'h25;
ROM_MEM[8102] = 8'hC1;
ROM_MEM[8103] = 8'h82;
ROM_MEM[8104] = 8'h09;
ROM_MEM[8105] = 8'h22;
ROM_MEM[8106] = 8'h80;
ROM_MEM[8107] = 8'h22;
ROM_MEM[8108] = 8'h81;
ROM_MEM[8109] = 8'h8E;
ROM_MEM[8110] = 8'h04;
ROM_MEM[8111] = 8'h26;
ROM_MEM[8112] = 8'h40;
ROM_MEM[8113] = 8'h8F;
ROM_MEM[8114] = 8'h00;
ROM_MEM[8115] = 8'h29;
ROM_MEM[8116] = 8'h80;
ROM_MEM[8117] = 8'h29;
ROM_MEM[8118] = 8'h81;
ROM_MEM[8119] = 8'h28;
ROM_MEM[8120] = 8'hC0;
ROM_MEM[8121] = 8'h28;
ROM_MEM[8122] = 8'h40;
ROM_MEM[8123] = 8'h26;
ROM_MEM[8124] = 8'hC0;
ROM_MEM[8125] = 8'h26;
ROM_MEM[8126] = 8'hC1;
ROM_MEM[8127] = 8'h26;
ROM_MEM[8128] = 8'hC1;
ROM_MEM[8129] = 8'h26;
ROM_MEM[8130] = 8'hC1;
ROM_MEM[8131] = 8'h26;
ROM_MEM[8132] = 8'hC1;
ROM_MEM[8133] = 8'h26;
ROM_MEM[8134] = 8'h41;
ROM_MEM[8135] = 8'h83;
ROM_MEM[8136] = 8'hFF;
ROM_MEM[8137] = 8'h26;
ROM_MEM[8138] = 8'h41;
ROM_MEM[8139] = 8'h83;
ROM_MEM[8140] = 8'hFF;
ROM_MEM[8141] = 8'h26;
ROM_MEM[8142] = 8'h41;
ROM_MEM[8143] = 8'h83;
ROM_MEM[8144] = 8'hFF;
ROM_MEM[8145] = 8'h26;
ROM_MEM[8146] = 8'h41;
ROM_MEM[8147] = 8'h00;
ROM_MEM[8148] = 8'h00;
ROM_MEM[8149] = 8'h80;
ROM_MEM[8150] = 8'h87;
ROM_MEM[8151] = 8'h87;
ROM_MEM[8152] = 8'h03;
ROM_MEM[8153] = 8'h42;
ROM_MEM[8154] = 8'hC0;
ROM_MEM[8155] = 8'h3F;
ROM_MEM[8156] = 8'h40;
ROM_MEM[8157] = 8'h00;
ROM_MEM[8158] = 8'h60;
ROM_MEM[8159] = 8'h42;
ROM_MEM[8160] = 8'h20;
ROM_MEM[8161] = 8'h42;
ROM_MEM[8162] = 8'hC0;
ROM_MEM[8163] = 8'h3F;
ROM_MEM[8164] = 8'h40;
ROM_MEM[8165] = 8'h00;
ROM_MEM[8166] = 8'h60;
ROM_MEM[8167] = 8'h45;
ROM_MEM[8168] = 8'h20;
ROM_MEM[8169] = 8'h45;
ROM_MEM[8170] = 8'hC0;
ROM_MEM[8171] = 8'h45;
ROM_MEM[8172] = 8'h61;
ROM_MEM[8173] = 8'h44;
ROM_MEM[8174] = 8'h40;
ROM_MEM[8175] = 8'h45;
ROM_MEM[8176] = 8'h10;
ROM_MEM[8177] = 8'h44;
ROM_MEM[8178] = 8'h10;
ROM_MEM[8179] = 8'h80;
ROM_MEM[8180] = 8'h5A;
ROM_MEM[8181] = 8'h42;
ROM_MEM[8182] = 8'h20;
ROM_MEM[8183] = 8'h3F;
ROM_MEM[8184] = 8'h60;
ROM_MEM[8185] = 8'h3F;
ROM_MEM[8186] = 8'h81;
ROM_MEM[8187] = 8'h3F;
ROM_MEM[8188] = 8'hC1;
ROM_MEM[8189] = 8'h00;
ROM_MEM[8190] = 8'h30;
ROM_MEM[8191] = 8'h42;
ROM_MEM[8192 ] = 8'h10;
ROM_MEM[8193 ] = 8'h42;
ROM_MEM[8194 ] = 8'h80;
ROM_MEM[8195 ] = 8'h3F;
ROM_MEM[8196 ] = 8'h40;
ROM_MEM[8197 ] = 8'h00;
ROM_MEM[8198 ] = 8'h30;
ROM_MEM[8199 ] = 8'h42;
ROM_MEM[8200 ] = 8'h10;
ROM_MEM[8201 ] = 8'h42;
ROM_MEM[8202 ] = 8'h80;
ROM_MEM[8203 ] = 8'h3F;
ROM_MEM[8204 ] = 8'h40;
ROM_MEM[8205 ] = 8'h00;
ROM_MEM[8206 ] = 8'h30;
ROM_MEM[8207 ] = 8'h45;
ROM_MEM[8208 ] = 8'h10;
ROM_MEM[8209 ] = 8'h45;
ROM_MEM[8210 ] = 8'h80;
ROM_MEM[8211 ] = 8'h45;
ROM_MEM[8212 ] = 8'h81;
ROM_MEM[8213 ] = 8'h45;
ROM_MEM[8214 ] = 8'hC1;
ROM_MEM[8215 ] = 8'h44;
ROM_MEM[8216 ] = 8'h20;
ROM_MEM[8217 ] = 8'h45;
ROM_MEM[8218 ] = 8'h10;
ROM_MEM[8219 ] = 8'h44;
ROM_MEM[8220 ] = 8'h10;
ROM_MEM[8221 ] = 8'h42;
ROM_MEM[8222 ] = 8'h20;
ROM_MEM[8223 ] = 8'h3F;
ROM_MEM[8224 ] = 8'h60;
ROM_MEM[8225 ] = 8'h83;
ROM_MEM[8226 ] = 8'hFF;
ROM_MEM[8227 ] = 8'h3F;
ROM_MEM[8228 ] = 8'h41;
ROM_MEM[8229 ] = 8'h83;
ROM_MEM[8230 ] = 8'hFF;
ROM_MEM[8231 ] = 8'h3F;
ROM_MEM[8232 ] = 8'h41;
ROM_MEM[8233 ] = 8'h83;
ROM_MEM[8234 ] = 8'hFF;
ROM_MEM[8235 ] = 8'h3F;
ROM_MEM[8236 ] = 8'h41;
ROM_MEM[8237 ] = 8'h83;
ROM_MEM[8238 ] = 8'hFF;
ROM_MEM[8239 ] = 8'h3F;
ROM_MEM[8240 ] = 8'h41;
ROM_MEM[8241 ] = 8'h83;
ROM_MEM[8242 ] = 8'hFF;
ROM_MEM[8243 ] = 8'h3F;
ROM_MEM[8244 ] = 8'h41;
ROM_MEM[8245 ] = 8'h00;
ROM_MEM[8246 ] = 8'h00;
ROM_MEM[8247 ] = 8'h80;
ROM_MEM[8248 ] = 8'h87;
ROM_MEM[8249 ] = 8'h87;
ROM_MEM[8250 ] = 8'h03;
ROM_MEM[8251 ] = 8'h3F;
ROM_MEM[8252 ] = 8'hC0;
ROM_MEM[8253 ] = 8'h3C;
ROM_MEM[8254 ] = 8'h40;
ROM_MEM[8255 ] = 8'h00;
ROM_MEM[8256 ] = 8'h60;
ROM_MEM[8257 ] = 8'h3F;
ROM_MEM[8258 ] = 8'h20;
ROM_MEM[8259 ] = 8'h3F;
ROM_MEM[8260 ] = 8'hC0;
ROM_MEM[8261 ] = 8'h3C;
ROM_MEM[8262 ] = 8'h40;
ROM_MEM[8263 ] = 8'h00;
ROM_MEM[8264 ] = 8'h60;
ROM_MEM[8265 ] = 8'h42;
ROM_MEM[8266 ] = 8'h20;
ROM_MEM[8267 ] = 8'h42;
ROM_MEM[8268 ] = 8'hC0;
ROM_MEM[8269 ] = 8'h42;
ROM_MEM[8270 ] = 8'h61;
ROM_MEM[8271 ] = 8'h41;
ROM_MEM[8272 ] = 8'h40;
ROM_MEM[8273 ] = 8'h42;
ROM_MEM[8274 ] = 8'h10;
ROM_MEM[8275 ] = 8'h41;
ROM_MEM[8276 ] = 8'h10;
ROM_MEM[8277 ] = 8'h80;
ROM_MEM[8278 ] = 8'h5A;
ROM_MEM[8279 ] = 8'h3F;
ROM_MEM[8280 ] = 8'h20;
ROM_MEM[8281 ] = 8'h3C;
ROM_MEM[8282 ] = 8'h60;
ROM_MEM[8283 ] = 8'h3C;
ROM_MEM[8284 ] = 8'h81;
ROM_MEM[8285 ] = 8'h3C;
ROM_MEM[8286 ] = 8'hC1;
ROM_MEM[8287 ] = 8'h00;
ROM_MEM[8288 ] = 8'h30;
ROM_MEM[8289 ] = 8'h3F;
ROM_MEM[8290 ] = 8'h10;
ROM_MEM[8291 ] = 8'h3F;
ROM_MEM[8292 ] = 8'h80;
ROM_MEM[8293 ] = 8'h3C;
ROM_MEM[8294 ] = 8'h40;
ROM_MEM[8295 ] = 8'h00;
ROM_MEM[8296 ] = 8'h30;
ROM_MEM[8297 ] = 8'h3F;
ROM_MEM[8298 ] = 8'h10;
ROM_MEM[8299 ] = 8'h3F;
ROM_MEM[8300 ] = 8'h80;
ROM_MEM[8301 ] = 8'h3C;
ROM_MEM[8302 ] = 8'h40;
ROM_MEM[8303 ] = 8'h00;
ROM_MEM[8304 ] = 8'h30;
ROM_MEM[8305 ] = 8'h42;
ROM_MEM[8306 ] = 8'h10;
ROM_MEM[8307 ] = 8'h42;
ROM_MEM[8308 ] = 8'h80;
ROM_MEM[8309 ] = 8'h42;
ROM_MEM[8310 ] = 8'h81;
ROM_MEM[8311 ] = 8'h42;
ROM_MEM[8312 ] = 8'hC1;
ROM_MEM[8313 ] = 8'h41;
ROM_MEM[8314 ] = 8'h20;
ROM_MEM[8315 ] = 8'h42;
ROM_MEM[8316 ] = 8'h10;
ROM_MEM[8317 ] = 8'h41;
ROM_MEM[8318 ] = 8'h10;
ROM_MEM[8319 ] = 8'h3F;
ROM_MEM[8320 ] = 8'h20;
ROM_MEM[8321 ] = 8'h3C;
ROM_MEM[8322 ] = 8'h60;
ROM_MEM[8323 ] = 8'h83;
ROM_MEM[8324 ] = 8'hFF;
ROM_MEM[8325 ] = 8'h3C;
ROM_MEM[8326 ] = 8'h41;
ROM_MEM[8327 ] = 8'h83;
ROM_MEM[8328 ] = 8'hFF;
ROM_MEM[8329 ] = 8'h3C;
ROM_MEM[8330 ] = 8'h41;
ROM_MEM[8331 ] = 8'h83;
ROM_MEM[8332 ] = 8'hFF;
ROM_MEM[8333 ] = 8'h3C;
ROM_MEM[8334 ] = 8'h41;
ROM_MEM[8335 ] = 8'h83;
ROM_MEM[8336 ] = 8'hFF;
ROM_MEM[8337 ] = 8'h3C;
ROM_MEM[8338 ] = 8'h41;
ROM_MEM[8339 ] = 8'h83;
ROM_MEM[8340 ] = 8'hFF;
ROM_MEM[8341 ] = 8'h3C;
ROM_MEM[8342 ] = 8'h41;
ROM_MEM[8343 ] = 8'h00;
ROM_MEM[8344 ] = 8'h00;
ROM_MEM[8345 ] = 8'h80;
ROM_MEM[8346 ] = 8'h87;
ROM_MEM[8347 ] = 8'h87;
ROM_MEM[8348 ] = 8'h03;
ROM_MEM[8349 ] = 8'h3B;
ROM_MEM[8350 ] = 8'hC0;
ROM_MEM[8351 ] = 8'h38;
ROM_MEM[8352 ] = 8'h40;
ROM_MEM[8353 ] = 8'h00;
ROM_MEM[8354 ] = 8'h60;
ROM_MEM[8355 ] = 8'h3B;
ROM_MEM[8356 ] = 8'h20;
ROM_MEM[8357 ] = 8'h3B;
ROM_MEM[8358 ] = 8'hC0;
ROM_MEM[8359 ] = 8'h38;
ROM_MEM[8360 ] = 8'h40;
ROM_MEM[8361 ] = 8'h00;
ROM_MEM[8362 ] = 8'h60;
ROM_MEM[8363 ] = 8'h3E;
ROM_MEM[8364 ] = 8'h20;
ROM_MEM[8365 ] = 8'h3E;
ROM_MEM[8366 ] = 8'hC0;
ROM_MEM[8367 ] = 8'h3E;
ROM_MEM[8368 ] = 8'h61;
ROM_MEM[8369 ] = 8'h3D;
ROM_MEM[8370 ] = 8'h40;
ROM_MEM[8371 ] = 8'h3E;
ROM_MEM[8372 ] = 8'h10;
ROM_MEM[8373 ] = 8'h3D;
ROM_MEM[8374 ] = 8'h10;
ROM_MEM[8375 ] = 8'h80;
ROM_MEM[8376 ] = 8'h5A;
ROM_MEM[8377 ] = 8'h3B;
ROM_MEM[8378 ] = 8'h20;
ROM_MEM[8379 ] = 8'h00;
ROM_MEM[8380 ] = 8'h20;
ROM_MEM[8381 ] = 8'h83;
ROM_MEM[8382 ] = 8'hFC;
ROM_MEM[8383 ] = 8'h8E;
ROM_MEM[8384 ] = 8'h02;
ROM_MEM[8385 ] = 8'h31;
ROM_MEM[8386 ] = 8'h10;
ROM_MEM[8387 ] = 8'h30;
ROM_MEM[8388 ] = 8'h10;
ROM_MEM[8389 ] = 8'h2E;
ROM_MEM[8390 ] = 8'h10;
ROM_MEM[8391 ] = 8'h2C;
ROM_MEM[8392 ] = 8'h10;
ROM_MEM[8393 ] = 8'h8F;
ROM_MEM[8394 ] = 8'h00;
ROM_MEM[8395 ] = 8'h36;
ROM_MEM[8396 ] = 8'h10;
ROM_MEM[8397 ] = 8'h35;
ROM_MEM[8398 ] = 8'h10;
ROM_MEM[8399 ] = 8'h33;
ROM_MEM[8400 ] = 8'h10;
ROM_MEM[8401 ] = 8'h31;
ROM_MEM[8402 ] = 8'h10;
ROM_MEM[8403 ] = 8'h8E;
ROM_MEM[8404 ] = 8'h03;
ROM_MEM[8405 ] = 8'h31;
ROM_MEM[8406 ] = 8'h10;
ROM_MEM[8407 ] = 8'h30;
ROM_MEM[8408 ] = 8'h10;
ROM_MEM[8409 ] = 8'h2E;
ROM_MEM[8410 ] = 8'h10;
ROM_MEM[8411 ] = 8'h2C;
ROM_MEM[8412 ] = 8'h10;
ROM_MEM[8413 ] = 8'h8F;
ROM_MEM[8414 ] = 8'h00;
ROM_MEM[8415 ] = 8'h36;
ROM_MEM[8416 ] = 8'h10;
ROM_MEM[8417 ] = 8'h35;
ROM_MEM[8418 ] = 8'h10;
ROM_MEM[8419 ] = 8'h33;
ROM_MEM[8420 ] = 8'h10;
ROM_MEM[8421 ] = 8'h31;
ROM_MEM[8422 ] = 8'h10;
ROM_MEM[8423 ] = 8'h83;
ROM_MEM[8424 ] = 8'h04;
ROM_MEM[8425 ] = 8'h3B;
ROM_MEM[8426 ] = 8'h80;
ROM_MEM[8427 ] = 8'h38;
ROM_MEM[8428 ] = 8'h40;
ROM_MEM[8429 ] = 8'h00;
ROM_MEM[8430 ] = 8'h30;
ROM_MEM[8431 ] = 8'h3B;
ROM_MEM[8432 ] = 8'h10;
ROM_MEM[8433 ] = 8'h3B;
ROM_MEM[8434 ] = 8'h80;
ROM_MEM[8435 ] = 8'h38;
ROM_MEM[8436 ] = 8'h40;
ROM_MEM[8437 ] = 8'h00;
ROM_MEM[8438 ] = 8'h40;
ROM_MEM[8439 ] = 8'h83;
ROM_MEM[8440 ] = 8'hFC;
ROM_MEM[8441 ] = 8'h00;
ROM_MEM[8442 ] = 8'h30;
ROM_MEM[8443 ] = 8'h2D;
ROM_MEM[8444 ] = 8'h10;
ROM_MEM[8445 ] = 8'h8E;
ROM_MEM[8446 ] = 8'h02;
ROM_MEM[8447 ] = 8'h32;
ROM_MEM[8448 ] = 8'h10;
ROM_MEM[8449 ] = 8'h31;
ROM_MEM[8450 ] = 8'h10;
ROM_MEM[8451 ] = 8'h2F;
ROM_MEM[8452 ] = 8'h10;
ROM_MEM[8453 ] = 8'h2D;
ROM_MEM[8454 ] = 8'h10;
ROM_MEM[8455 ] = 8'h32;
ROM_MEM[8456 ] = 8'h10;
ROM_MEM[8457 ] = 8'h31;
ROM_MEM[8458 ] = 8'h10;
ROM_MEM[8459 ] = 8'h2F;
ROM_MEM[8460 ] = 8'h10;
ROM_MEM[8461 ] = 8'h2D;
ROM_MEM[8462 ] = 8'h10;
ROM_MEM[8463 ] = 8'h39;
ROM_MEM[8464 ] = 8'h10;
ROM_MEM[8465 ] = 8'h38;
ROM_MEM[8466 ] = 8'h10;
ROM_MEM[8467 ] = 8'h36;
ROM_MEM[8468 ] = 8'h10;
ROM_MEM[8469 ] = 8'h34;
ROM_MEM[8470 ] = 8'h10;
ROM_MEM[8471 ] = 8'h8F;
ROM_MEM[8472 ] = 8'h00;
ROM_MEM[8473 ] = 8'h38;
ROM_MEM[8474 ] = 8'h20;
ROM_MEM[8475 ] = 8'h00;
ROM_MEM[8476 ] = 8'h20;
ROM_MEM[8477 ] = 8'h00;
ROM_MEM[8478 ] = 8'h40;
ROM_MEM[8479 ] = 8'h83;
ROM_MEM[8480 ] = 8'hFF;
ROM_MEM[8481 ] = 8'h8E;
ROM_MEM[8482 ] = 8'h02;
ROM_MEM[8483 ] = 8'h38;
ROM_MEM[8484 ] = 8'h10;
ROM_MEM[8485 ] = 8'h36;
ROM_MEM[8486 ] = 8'h10;
ROM_MEM[8487 ] = 8'h35;
ROM_MEM[8488 ] = 8'h10;
ROM_MEM[8489 ] = 8'h33;
ROM_MEM[8490 ] = 8'h10;
ROM_MEM[8491 ] = 8'h8F;
ROM_MEM[8492 ] = 8'h00;
ROM_MEM[8493 ] = 8'h83;
ROM_MEM[8494 ] = 8'hFF;
ROM_MEM[8495 ] = 8'h8E;
ROM_MEM[8496 ] = 8'h03;
ROM_MEM[8497 ] = 8'h86;
ROM_MEM[8498 ] = 8'h01;
ROM_MEM[8499 ] = 8'h3F;
ROM_MEM[8500 ] = 8'h10;
ROM_MEM[8501 ] = 8'h86;
ROM_MEM[8502 ] = 8'h00;
ROM_MEM[8503 ] = 8'h3D;
ROM_MEM[8504 ] = 8'h10;
ROM_MEM[8505 ] = 8'h86;
ROM_MEM[8506 ] = 8'h01;
ROM_MEM[8507 ] = 8'h3C;
ROM_MEM[8508 ] = 8'h10;
ROM_MEM[8509 ] = 8'h86;
ROM_MEM[8510 ] = 8'h00;
ROM_MEM[8511 ] = 8'h3A;
ROM_MEM[8512 ] = 8'h10;
ROM_MEM[8513 ] = 8'h8F;
ROM_MEM[8514 ] = 8'h00;
ROM_MEM[8515 ] = 8'h38;
ROM_MEM[8516 ] = 8'h20;
ROM_MEM[8517 ] = 8'h00;
ROM_MEM[8518 ] = 8'h20;
ROM_MEM[8519 ] = 8'h00;
ROM_MEM[8520 ] = 8'h00;
ROM_MEM[8521 ] = 8'h80;
ROM_MEM[8522 ] = 8'h87;
ROM_MEM[8523 ] = 8'h87;
ROM_MEM[8524 ] = 8'h03;
ROM_MEM[8525 ] = 8'h00;
ROM_MEM[8526 ] = 8'h60;
ROM_MEM[8527 ] = 8'h20;
ROM_MEM[8528 ] = 8'hC0;
ROM_MEM[8529 ] = 8'h20;
ROM_MEM[8530 ] = 8'h60;
ROM_MEM[8531 ] = 8'h20;
ROM_MEM[8532 ] = 8'h61;
ROM_MEM[8533 ] = 8'h20;
ROM_MEM[8534 ] = 8'hC0;
ROM_MEM[8535 ] = 8'h20;
ROM_MEM[8536 ] = 8'h60;
ROM_MEM[8537 ] = 8'h20;
ROM_MEM[8538 ] = 8'h21;
ROM_MEM[8539 ] = 8'h00;
ROM_MEM[8540 ] = 8'h40;
ROM_MEM[8541 ] = 8'h20;
ROM_MEM[8542 ] = 8'h20;
ROM_MEM[8543 ] = 8'h00;
ROM_MEM[8544 ] = 8'h40;
ROM_MEM[8545 ] = 8'h20;
ROM_MEM[8546 ] = 8'h20;
ROM_MEM[8547 ] = 8'h00;
ROM_MEM[8548 ] = 8'h40;
ROM_MEM[8549 ] = 8'h20;
ROM_MEM[8550 ] = 8'h20;
ROM_MEM[8551 ] = 8'h00;
ROM_MEM[8552 ] = 8'h40;
ROM_MEM[8553 ] = 8'h80;
ROM_MEM[8554 ] = 8'h5A;
ROM_MEM[8555 ] = 8'h25;
ROM_MEM[8556 ] = 8'h20;
ROM_MEM[8557 ] = 8'h00;
ROM_MEM[8558 ] = 8'h20;
ROM_MEM[8559 ] = 8'h25;
ROM_MEM[8560 ] = 8'h40;
ROM_MEM[8561 ] = 8'h25;
ROM_MEM[8562 ] = 8'h40;
ROM_MEM[8563 ] = 8'h25;
ROM_MEM[8564 ] = 8'h40;
ROM_MEM[8565 ] = 8'h8E;
ROM_MEM[8566 ] = 8'h06;
ROM_MEM[8567 ] = 8'h25;
ROM_MEM[8568 ] = 8'h40;
ROM_MEM[8569 ] = 8'h25;
ROM_MEM[8570 ] = 8'h40;
ROM_MEM[8571 ] = 8'h25;
ROM_MEM[8572 ] = 8'h40;
ROM_MEM[8573 ] = 8'h25;
ROM_MEM[8574 ] = 8'h40;
ROM_MEM[8575 ] = 8'h8F;
ROM_MEM[8576 ] = 8'h00;
ROM_MEM[8577 ] = 8'h8E;
ROM_MEM[8578 ] = 8'h03;
ROM_MEM[8579 ] = 8'h83;
ROM_MEM[8580 ] = 8'hFF;
ROM_MEM[8581 ] = 8'h25;
ROM_MEM[8582 ] = 8'h40;
ROM_MEM[8583 ] = 8'h8F;
ROM_MEM[8584 ] = 8'h00;
ROM_MEM[8585 ] = 8'h00;
ROM_MEM[8586 ] = 8'h00;
ROM_MEM[8587 ] = 8'h80;
ROM_MEM[8588 ] = 8'h98;
ROM_MEM[8589 ] = 8'h87;
ROM_MEM[8590 ] = 8'h03;
ROM_MEM[8591 ] = 8'h42;
ROM_MEM[8592 ] = 8'h16;
ROM_MEM[8593 ] = 8'h8E;
ROM_MEM[8594 ] = 8'h02;
ROM_MEM[8595 ] = 8'h42;
ROM_MEM[8596 ] = 8'h80;
ROM_MEM[8597 ] = 8'h3F;
ROM_MEM[8598 ] = 8'h20;
ROM_MEM[8599 ] = 8'h00;
ROM_MEM[8600 ] = 8'h20;
ROM_MEM[8601 ] = 8'h3F;
ROM_MEM[8602 ] = 8'h16;
ROM_MEM[8603 ] = 8'h3F;
ROM_MEM[8604 ] = 8'h16;
ROM_MEM[8605 ] = 8'h3F;
ROM_MEM[8606 ] = 8'h14;
ROM_MEM[8607 ] = 8'h8F;
ROM_MEM[8608 ] = 8'h00;
ROM_MEM[8609 ] = 8'h45;
ROM_MEM[8610 ] = 8'h80;
ROM_MEM[8611 ] = 8'h44;
ROM_MEM[8612 ] = 8'h40;
ROM_MEM[8613 ] = 8'h44;
ROM_MEM[8614 ] = 8'h16;
ROM_MEM[8615 ] = 8'h45;
ROM_MEM[8616 ] = 8'h16;
ROM_MEM[8617 ] = 8'h44;
ROM_MEM[8618 ] = 8'h14;
ROM_MEM[8619 ] = 8'h42;
ROM_MEM[8620 ] = 8'h40;
ROM_MEM[8621 ] = 8'h3F;
ROM_MEM[8622 ] = 8'hC0;
ROM_MEM[8623 ] = 8'h3F;
ROM_MEM[8624 ] = 8'h81;
ROM_MEM[8625 ] = 8'h3F;
ROM_MEM[8626 ] = 8'h21;
ROM_MEM[8627 ] = 8'h00;
ROM_MEM[8628 ] = 8'h20;
ROM_MEM[8629 ] = 8'h00;
ROM_MEM[8630 ] = 8'h16;
ROM_MEM[8631 ] = 8'h00;
ROM_MEM[8632 ] = 8'h16;
ROM_MEM[8633 ] = 8'h42;
ROM_MEM[8634 ] = 8'h14;
ROM_MEM[8635 ] = 8'h8E;
ROM_MEM[8636 ] = 8'h02;
ROM_MEM[8637 ] = 8'h42;
ROM_MEM[8638 ] = 8'h80;
ROM_MEM[8639 ] = 8'h3F;
ROM_MEM[8640 ] = 8'h20;
ROM_MEM[8641 ] = 8'h00;
ROM_MEM[8642 ] = 8'h20;
ROM_MEM[8643 ] = 8'h3F;
ROM_MEM[8644 ] = 8'h16;
ROM_MEM[8645 ] = 8'h3F;
ROM_MEM[8646 ] = 8'h16;
ROM_MEM[8647 ] = 8'h3F;
ROM_MEM[8648 ] = 8'h14;
ROM_MEM[8649 ] = 8'h8F;
ROM_MEM[8650 ] = 8'h00;
ROM_MEM[8651 ] = 8'h45;
ROM_MEM[8652 ] = 8'h80;
ROM_MEM[8653 ] = 8'h44;
ROM_MEM[8654 ] = 8'h20;
ROM_MEM[8655 ] = 8'h00;
ROM_MEM[8656 ] = 8'h20;
ROM_MEM[8657 ] = 8'h44;
ROM_MEM[8658 ] = 8'h16;
ROM_MEM[8659 ] = 8'h45;
ROM_MEM[8660 ] = 8'h16;
ROM_MEM[8661 ] = 8'h44;
ROM_MEM[8662 ] = 8'h14;
ROM_MEM[8663 ] = 8'h8E;
ROM_MEM[8664 ] = 8'h02;
ROM_MEM[8665 ] = 8'h42;
ROM_MEM[8666 ] = 8'h40;
ROM_MEM[8667 ] = 8'h3F;
ROM_MEM[8668 ] = 8'h40;
ROM_MEM[8669 ] = 8'h45;
ROM_MEM[8670 ] = 8'h40;
ROM_MEM[8671 ] = 8'h44;
ROM_MEM[8672 ] = 8'h16;
ROM_MEM[8673 ] = 8'h45;
ROM_MEM[8674 ] = 8'h16;
ROM_MEM[8675 ] = 8'h44;
ROM_MEM[8676 ] = 8'h14;
ROM_MEM[8677 ] = 8'h8F;
ROM_MEM[8678 ] = 8'h00;
ROM_MEM[8679 ] = 8'h8E;
ROM_MEM[8680 ] = 8'h02;
ROM_MEM[8681 ] = 8'h42;
ROM_MEM[8682 ] = 8'h40;
ROM_MEM[8683 ] = 8'h44;
ROM_MEM[8684 ] = 8'h16;
ROM_MEM[8685 ] = 8'h45;
ROM_MEM[8686 ] = 8'h16;
ROM_MEM[8687 ] = 8'h44;
ROM_MEM[8688 ] = 8'h14;
ROM_MEM[8689 ] = 8'h8F;
ROM_MEM[8690 ] = 8'h00;
ROM_MEM[8691 ] = 8'h42;
ROM_MEM[8692 ] = 8'h40;
ROM_MEM[8693 ] = 8'h45;
ROM_MEM[8694 ] = 8'h16;
ROM_MEM[8695 ] = 8'h44;
ROM_MEM[8696 ] = 8'h16;
ROM_MEM[8697 ] = 8'h45;
ROM_MEM[8698 ] = 8'h14;
ROM_MEM[8699 ] = 8'h46;
ROM_MEM[8700 ] = 8'h80;
ROM_MEM[8701 ] = 8'h46;
ROM_MEM[8702 ] = 8'h81;
ROM_MEM[8703 ] = 8'h46;
ROM_MEM[8704 ] = 8'hC1;
ROM_MEM[8705 ] = 8'h00;
ROM_MEM[8706 ] = 8'h00;
ROM_MEM[8707 ] = 8'h80;
ROM_MEM[8708 ] = 8'h98;
ROM_MEM[8709 ] = 8'h87;
ROM_MEM[8710 ] = 8'h03;
ROM_MEM[8711 ] = 8'h3F;
ROM_MEM[8712 ] = 8'h16;
ROM_MEM[8713 ] = 8'h8E;
ROM_MEM[8714 ] = 8'h02;
ROM_MEM[8715 ] = 8'h3F;
ROM_MEM[8716 ] = 8'h80;
ROM_MEM[8717 ] = 8'h3C;
ROM_MEM[8718 ] = 8'h20;
ROM_MEM[8719 ] = 8'h00;
ROM_MEM[8720 ] = 8'h20;
ROM_MEM[8721 ] = 8'h3C;
ROM_MEM[8722 ] = 8'h16;
ROM_MEM[8723 ] = 8'h3C;
ROM_MEM[8724 ] = 8'h16;
ROM_MEM[8725 ] = 8'h3C;
ROM_MEM[8726 ] = 8'h14;
ROM_MEM[8727 ] = 8'h8F;
ROM_MEM[8728 ] = 8'h00;
ROM_MEM[8729 ] = 8'h42;
ROM_MEM[8730 ] = 8'h80;
ROM_MEM[8731 ] = 8'h41;
ROM_MEM[8732 ] = 8'h40;
ROM_MEM[8733 ] = 8'h41;
ROM_MEM[8734 ] = 8'h16;
ROM_MEM[8735 ] = 8'h42;
ROM_MEM[8736 ] = 8'h16;
ROM_MEM[8737 ] = 8'h41;
ROM_MEM[8738 ] = 8'h14;
ROM_MEM[8739 ] = 8'h3F;
ROM_MEM[8740 ] = 8'h40;
ROM_MEM[8741 ] = 8'h3C;
ROM_MEM[8742 ] = 8'hC0;
ROM_MEM[8743 ] = 8'h3C;
ROM_MEM[8744 ] = 8'h81;
ROM_MEM[8745 ] = 8'h3C;
ROM_MEM[8746 ] = 8'h21;
ROM_MEM[8747 ] = 8'h00;
ROM_MEM[8748 ] = 8'h20;
ROM_MEM[8749 ] = 8'h00;
ROM_MEM[8750 ] = 8'h16;
ROM_MEM[8751 ] = 8'h00;
ROM_MEM[8752 ] = 8'h16;
ROM_MEM[8753 ] = 8'h3E;
ROM_MEM[8754 ] = 8'h14;
ROM_MEM[8755 ] = 8'h8E;
ROM_MEM[8756 ] = 8'h02;
ROM_MEM[8757 ] = 8'h3E;
ROM_MEM[8758 ] = 8'h80;
ROM_MEM[8759 ] = 8'h3B;
ROM_MEM[8760 ] = 8'h20;
ROM_MEM[8761 ] = 8'h00;
ROM_MEM[8762 ] = 8'h20;
ROM_MEM[8763 ] = 8'h3B;
ROM_MEM[8764 ] = 8'h16;
ROM_MEM[8765 ] = 8'h3B;
ROM_MEM[8766 ] = 8'h16;
ROM_MEM[8767 ] = 8'h3B;
ROM_MEM[8768 ] = 8'h14;
ROM_MEM[8769 ] = 8'h8F;
ROM_MEM[8770 ] = 8'h00;
ROM_MEM[8771 ] = 8'h42;
ROM_MEM[8772 ] = 8'h80;
ROM_MEM[8773 ] = 8'h41;
ROM_MEM[8774 ] = 8'h20;
ROM_MEM[8775 ] = 8'h00;
ROM_MEM[8776 ] = 8'h20;
ROM_MEM[8777 ] = 8'h41;
ROM_MEM[8778 ] = 8'h16;
ROM_MEM[8779 ] = 8'h42;
ROM_MEM[8780 ] = 8'h16;
ROM_MEM[8781 ] = 8'h41;
ROM_MEM[8782 ] = 8'h14;
ROM_MEM[8783 ] = 8'h8E;
ROM_MEM[8784 ] = 8'h02;
ROM_MEM[8785 ] = 8'h3F;
ROM_MEM[8786 ] = 8'h40;
ROM_MEM[8787 ] = 8'h3C;
ROM_MEM[8788 ] = 8'h40;
ROM_MEM[8789 ] = 8'h42;
ROM_MEM[8790 ] = 8'h40;
ROM_MEM[8791 ] = 8'h41;
ROM_MEM[8792 ] = 8'h16;
ROM_MEM[8793 ] = 8'h42;
ROM_MEM[8794 ] = 8'h16;
ROM_MEM[8795 ] = 8'h41;
ROM_MEM[8796 ] = 8'h14;
ROM_MEM[8797 ] = 8'h8F;
ROM_MEM[8798 ] = 8'h00;
ROM_MEM[8799 ] = 8'h8E;
ROM_MEM[8800 ] = 8'h02;
ROM_MEM[8801 ] = 8'h3E;
ROM_MEM[8802 ] = 8'h40;
ROM_MEM[8803 ] = 8'h41;
ROM_MEM[8804 ] = 8'h16;
ROM_MEM[8805 ] = 8'h42;
ROM_MEM[8806 ] = 8'h16;
ROM_MEM[8807 ] = 8'h41;
ROM_MEM[8808 ] = 8'h14;
ROM_MEM[8809 ] = 8'h8F;
ROM_MEM[8810 ] = 8'h00;
ROM_MEM[8811 ] = 8'h3E;
ROM_MEM[8812 ] = 8'h40;
ROM_MEM[8813 ] = 8'h42;
ROM_MEM[8814 ] = 8'h16;
ROM_MEM[8815 ] = 8'h41;
ROM_MEM[8816 ] = 8'h16;
ROM_MEM[8817 ] = 8'h42;
ROM_MEM[8818 ] = 8'h14;
ROM_MEM[8819 ] = 8'h43;
ROM_MEM[8820 ] = 8'h80;
ROM_MEM[8821 ] = 8'h43;
ROM_MEM[8822 ] = 8'h81;
ROM_MEM[8823 ] = 8'h43;
ROM_MEM[8824 ] = 8'hC1;
ROM_MEM[8825 ] = 8'h00;
ROM_MEM[8826 ] = 8'h00;
ROM_MEM[8827 ] = 8'h80;
ROM_MEM[8828 ] = 8'h98;
ROM_MEM[8829 ] = 8'h87;
ROM_MEM[8830 ] = 8'h03;
ROM_MEM[8831 ] = 8'h3B;
ROM_MEM[8832 ] = 8'h16;
ROM_MEM[8833 ] = 8'h8E;
ROM_MEM[8834 ] = 8'h02;
ROM_MEM[8835 ] = 8'h3B;
ROM_MEM[8836 ] = 8'h80;
ROM_MEM[8837 ] = 8'h38;
ROM_MEM[8838 ] = 8'h20;
ROM_MEM[8839 ] = 8'h00;
ROM_MEM[8840 ] = 8'h20;
ROM_MEM[8841 ] = 8'h38;
ROM_MEM[8842 ] = 8'h16;
ROM_MEM[8843 ] = 8'h38;
ROM_MEM[8844 ] = 8'h16;
ROM_MEM[8845 ] = 8'h38;
ROM_MEM[8846 ] = 8'h14;
ROM_MEM[8847 ] = 8'h8F;
ROM_MEM[8848 ] = 8'h00;
ROM_MEM[8849 ] = 8'h3E;
ROM_MEM[8850 ] = 8'h80;
ROM_MEM[8851 ] = 8'h3D;
ROM_MEM[8852 ] = 8'h40;
ROM_MEM[8853 ] = 8'h3D;
ROM_MEM[8854 ] = 8'h16;
ROM_MEM[8855 ] = 8'h3E;
ROM_MEM[8856 ] = 8'h16;
ROM_MEM[8857 ] = 8'h3D;
ROM_MEM[8858 ] = 8'h14;
ROM_MEM[8859 ] = 8'h3B;
ROM_MEM[8860 ] = 8'h40;
ROM_MEM[8861 ] = 8'h38;
ROM_MEM[8862 ] = 8'hC0;
ROM_MEM[8863 ] = 8'h38;
ROM_MEM[8864 ] = 8'h81;
ROM_MEM[8865 ] = 8'h38;
ROM_MEM[8866 ] = 8'h21;
ROM_MEM[8867 ] = 8'h00;
ROM_MEM[8868 ] = 8'h20;
ROM_MEM[8869 ] = 8'h00;
ROM_MEM[8870 ] = 8'h16;
ROM_MEM[8871 ] = 8'h00;
ROM_MEM[8872 ] = 8'h16;
ROM_MEM[8873 ] = 8'h39;
ROM_MEM[8874 ] = 8'h14;
ROM_MEM[8875 ] = 8'h8E;
ROM_MEM[8876 ] = 8'h02;
ROM_MEM[8877 ] = 8'h39;
ROM_MEM[8878 ] = 8'h80;
ROM_MEM[8879 ] = 8'h36;
ROM_MEM[8880 ] = 8'h20;
ROM_MEM[8881 ] = 8'h00;
ROM_MEM[8882 ] = 8'h20;
ROM_MEM[8883 ] = 8'h36;
ROM_MEM[8884 ] = 8'h16;
ROM_MEM[8885 ] = 8'h36;
ROM_MEM[8886 ] = 8'h16;
ROM_MEM[8887 ] = 8'h36;
ROM_MEM[8888 ] = 8'h14;
ROM_MEM[8889 ] = 8'h8F;
ROM_MEM[8890 ] = 8'h00;
ROM_MEM[8891 ] = 8'h3E;
ROM_MEM[8892 ] = 8'h80;
ROM_MEM[8893 ] = 8'h3D;
ROM_MEM[8894 ] = 8'h20;
ROM_MEM[8895 ] = 8'h00;
ROM_MEM[8896 ] = 8'h20;
ROM_MEM[8897 ] = 8'h3D;
ROM_MEM[8898 ] = 8'h16;
ROM_MEM[8899 ] = 8'h3E;
ROM_MEM[8900 ] = 8'h16;
ROM_MEM[8901 ] = 8'h3D;
ROM_MEM[8902 ] = 8'h14;
ROM_MEM[8903 ] = 8'h8E;
ROM_MEM[8904 ] = 8'h02;
ROM_MEM[8905 ] = 8'h3B;
ROM_MEM[8906 ] = 8'h40;
ROM_MEM[8907 ] = 8'h38;
ROM_MEM[8908 ] = 8'h40;
ROM_MEM[8909 ] = 8'h3E;
ROM_MEM[8910 ] = 8'h40;
ROM_MEM[8911 ] = 8'h3D;
ROM_MEM[8912 ] = 8'h16;
ROM_MEM[8913 ] = 8'h3E;
ROM_MEM[8914 ] = 8'h16;
ROM_MEM[8915 ] = 8'h3D;
ROM_MEM[8916 ] = 8'h14;
ROM_MEM[8917 ] = 8'h8F;
ROM_MEM[8918 ] = 8'h00;
ROM_MEM[8919 ] = 8'h8E;
ROM_MEM[8920 ] = 8'h02;
ROM_MEM[8921 ] = 8'h39;
ROM_MEM[8922 ] = 8'h40;
ROM_MEM[8923 ] = 8'h3D;
ROM_MEM[8924 ] = 8'h16;
ROM_MEM[8925 ] = 8'h3E;
ROM_MEM[8926 ] = 8'h16;
ROM_MEM[8927 ] = 8'h3D;
ROM_MEM[8928 ] = 8'h14;
ROM_MEM[8929 ] = 8'h8F;
ROM_MEM[8930 ] = 8'h00;
ROM_MEM[8931 ] = 8'h39;
ROM_MEM[8932 ] = 8'h40;
ROM_MEM[8933 ] = 8'h3E;
ROM_MEM[8934 ] = 8'h16;
ROM_MEM[8935 ] = 8'h3D;
ROM_MEM[8936 ] = 8'h16;
ROM_MEM[8937 ] = 8'h3E;
ROM_MEM[8938 ] = 8'h14;
ROM_MEM[8939 ] = 8'h3F;
ROM_MEM[8940 ] = 8'h80;
ROM_MEM[8941 ] = 8'h3F;
ROM_MEM[8942 ] = 8'h81;
ROM_MEM[8943 ] = 8'h3F;
ROM_MEM[8944 ] = 8'hC1;
ROM_MEM[8945 ] = 8'h00;
ROM_MEM[8946 ] = 8'h00;
ROM_MEM[8947 ] = 8'h80;
ROM_MEM[8948 ] = 8'h98;
ROM_MEM[8949 ] = 8'h87;
ROM_MEM[8950 ] = 8'h02;
ROM_MEM[8951 ] = 8'h83;
ROM_MEM[8952 ] = 8'hFF;
ROM_MEM[8953 ] = 8'h00;
ROM_MEM[8954 ] = 8'h16;
ROM_MEM[8955 ] = 8'h8E;
ROM_MEM[8956 ] = 8'h0D;
ROM_MEM[8957 ] = 8'h25;
ROM_MEM[8958 ] = 8'h80;
ROM_MEM[8959 ] = 8'h25;
ROM_MEM[8960 ] = 8'h80;
ROM_MEM[8961 ] = 8'h8F;
ROM_MEM[8962 ] = 8'h00;
ROM_MEM[8963 ] = 8'h25;
ROM_MEM[8964 ] = 8'h40;
ROM_MEM[8965 ] = 8'h00;
ROM_MEM[8966 ] = 8'h00;
ROM_MEM[8967 ] = 8'h80;
ROM_MEM[8968 ] = 8'h5A;
ROM_MEM[8969 ] = 8'h87;
ROM_MEM[8970 ] = 8'h01;
ROM_MEM[8971 ] = 8'h33;
ROM_MEM[8972 ] = 8'h16;
ROM_MEM[8973 ] = 8'h33;
ROM_MEM[8974 ] = 8'h16;
ROM_MEM[8975 ] = 8'h33;
ROM_MEM[8976 ] = 8'h14;
ROM_MEM[8977 ] = 8'h87;
ROM_MEM[8978 ] = 8'h02;
ROM_MEM[8979 ] = 8'h38;
ROM_MEM[8980 ] = 8'h80;
ROM_MEM[8981 ] = 8'h3F;
ROM_MEM[8982 ] = 8'h80;
ROM_MEM[8983 ] = 8'h3D;
ROM_MEM[8984 ] = 8'h16;
ROM_MEM[8985 ] = 8'h3C;
ROM_MEM[8986 ] = 8'h16;
ROM_MEM[8987 ] = 8'h3A;
ROM_MEM[8988 ] = 8'h14;
ROM_MEM[8989 ] = 8'h44;
ROM_MEM[8990 ] = 8'h80;
ROM_MEM[8991 ] = 8'h3F;
ROM_MEM[8992 ] = 8'h40;
ROM_MEM[8993 ] = 8'h3D;
ROM_MEM[8994 ] = 8'h16;
ROM_MEM[8995 ] = 8'h3C;
ROM_MEM[8996 ] = 8'h16;
ROM_MEM[8997 ] = 8'h3A;
ROM_MEM[8998 ] = 8'h14;
ROM_MEM[8999 ] = 8'h44;
ROM_MEM[9000 ] = 8'h80;
ROM_MEM[9001 ] = 8'h3F;
ROM_MEM[9002 ] = 8'h40;
ROM_MEM[9003 ] = 8'h3D;
ROM_MEM[9004 ] = 8'h16;
ROM_MEM[9005 ] = 8'h3C;
ROM_MEM[9006 ] = 8'h16;
ROM_MEM[9007 ] = 8'h3D;
ROM_MEM[9008 ] = 8'h14;
ROM_MEM[9009 ] = 8'h3A;
ROM_MEM[9010 ] = 8'hC0;
ROM_MEM[9011 ] = 8'h00;
ROM_MEM[9012 ] = 8'h00;
ROM_MEM[9013 ] = 8'h80;
ROM_MEM[9014 ] = 8'h5A;
ROM_MEM[9015 ] = 8'h87;
ROM_MEM[9016 ] = 8'h01;
ROM_MEM[9017 ] = 8'h27;
ROM_MEM[9018 ] = 8'h16;
ROM_MEM[9019 ] = 8'h27;
ROM_MEM[9020 ] = 8'h16;
ROM_MEM[9021 ] = 8'h27;
ROM_MEM[9022 ] = 8'h14;
ROM_MEM[9023 ] = 8'h87;
ROM_MEM[9024 ] = 8'h02;
ROM_MEM[9025 ] = 8'h33;
ROM_MEM[9026 ] = 8'h80;
ROM_MEM[9027 ] = 8'h3C;
ROM_MEM[9028 ] = 8'h80;
ROM_MEM[9029 ] = 8'h38;
ROM_MEM[9030 ] = 8'h16;
ROM_MEM[9031 ] = 8'h00;
ROM_MEM[9032 ] = 8'h16;
ROM_MEM[9033 ] = 8'h00;
ROM_MEM[9034 ] = 8'h14;
ROM_MEM[9035 ] = 8'h3F;
ROM_MEM[9036 ] = 8'h80;
ROM_MEM[9037 ] = 8'h3C;
ROM_MEM[9038 ] = 8'h40;
ROM_MEM[9039 ] = 8'h38;
ROM_MEM[9040 ] = 8'h16;
ROM_MEM[9041 ] = 8'h00;
ROM_MEM[9042 ] = 8'h16;
ROM_MEM[9043 ] = 8'h00;
ROM_MEM[9044 ] = 8'h14;
ROM_MEM[9045 ] = 8'h3F;
ROM_MEM[9046 ] = 8'h80;
ROM_MEM[9047 ] = 8'h3C;
ROM_MEM[9048 ] = 8'h40;
ROM_MEM[9049 ] = 8'h3A;
ROM_MEM[9050 ] = 8'h16;
ROM_MEM[9051 ] = 8'h39;
ROM_MEM[9052 ] = 8'h16;
ROM_MEM[9053 ] = 8'h3A;
ROM_MEM[9054 ] = 8'h14;
ROM_MEM[9055 ] = 8'h37;
ROM_MEM[9056 ] = 8'hC0;
ROM_MEM[9057 ] = 8'h00;
ROM_MEM[9058 ] = 8'h00;
ROM_MEM[9059 ] = 8'h80;
ROM_MEM[9060 ] = 8'h5A;
ROM_MEM[9061 ] = 8'h87;
ROM_MEM[9062 ] = 8'h02;
ROM_MEM[9063 ] = 8'h00;
ROM_MEM[9064 ] = 8'h40;
ROM_MEM[9065 ] = 8'h30;
ROM_MEM[9066 ] = 8'h80;
ROM_MEM[9067 ] = 8'h38;
ROM_MEM[9068 ] = 8'h80;
ROM_MEM[9069 ] = 8'h35;
ROM_MEM[9070 ] = 8'h16;
ROM_MEM[9071 ] = 8'h00;
ROM_MEM[9072 ] = 8'h16;
ROM_MEM[9073 ] = 8'h00;
ROM_MEM[9074 ] = 8'h14;
ROM_MEM[9075 ] = 8'h3C;
ROM_MEM[9076 ] = 8'h80;
ROM_MEM[9077 ] = 8'h38;
ROM_MEM[9078 ] = 8'h40;
ROM_MEM[9079 ] = 8'h35;
ROM_MEM[9080 ] = 8'h16;
ROM_MEM[9081 ] = 8'h00;
ROM_MEM[9082 ] = 8'h16;
ROM_MEM[9083 ] = 8'h00;
ROM_MEM[9084 ] = 8'h14;
ROM_MEM[9085 ] = 8'h3C;
ROM_MEM[9086 ] = 8'h80;
ROM_MEM[9087 ] = 8'h38;
ROM_MEM[9088 ] = 8'h40;
ROM_MEM[9089 ] = 8'h36;
ROM_MEM[9090 ] = 8'h16;
ROM_MEM[9091 ] = 8'h35;
ROM_MEM[9092 ] = 8'h16;
ROM_MEM[9093 ] = 8'h36;
ROM_MEM[9094 ] = 8'h14;
ROM_MEM[9095 ] = 8'h00;
ROM_MEM[9096 ] = 8'h40;
ROM_MEM[9097 ] = 8'h27;
ROM_MEM[9098 ] = 8'h80;
ROM_MEM[9099 ] = 8'h00;
ROM_MEM[9100 ] = 8'h00;
ROM_MEM[9101 ] = 8'h80;
ROM_MEM[9102 ] = 8'h5A;
ROM_MEM[9103 ] = 8'h87;
ROM_MEM[9104 ] = 8'h01;
ROM_MEM[9105 ] = 8'h27;
ROM_MEM[9106 ] = 8'h16;
ROM_MEM[9107 ] = 8'h27;
ROM_MEM[9108 ] = 8'h16;
ROM_MEM[9109 ] = 8'h27;
ROM_MEM[9110 ] = 8'h14;
ROM_MEM[9111 ] = 8'h87;
ROM_MEM[9112 ] = 8'h02;
ROM_MEM[9113 ] = 8'h20;
ROM_MEM[9114 ] = 8'h40;
ROM_MEM[9115 ] = 8'h1F;
ROM_MEM[9116 ] = 8'h40;
ROM_MEM[9117 ] = 8'h1D;
ROM_MEM[9118 ] = 8'h40;
ROM_MEM[9119 ] = 8'h1B;
ROM_MEM[9120 ] = 8'h40;
ROM_MEM[9121 ] = 8'h19;
ROM_MEM[9122 ] = 8'h40;
ROM_MEM[9123 ] = 8'h20;
ROM_MEM[9124 ] = 8'h40;
ROM_MEM[9125 ] = 8'h1F;
ROM_MEM[9126 ] = 8'h40;
ROM_MEM[9127 ] = 8'h1D;
ROM_MEM[9128 ] = 8'h40;
ROM_MEM[9129 ] = 8'h1B;
ROM_MEM[9130 ] = 8'h40;
ROM_MEM[9131 ] = 8'h20;
ROM_MEM[9132 ] = 8'h40;
ROM_MEM[9133 ] = 8'h1F;
ROM_MEM[9134 ] = 8'h40;
ROM_MEM[9135 ] = 8'h1D;
ROM_MEM[9136 ] = 8'h40;
ROM_MEM[9137 ] = 8'h1E;
ROM_MEM[9138 ] = 8'h40;
ROM_MEM[9139 ] = 8'h1B;
ROM_MEM[9140 ] = 8'h40;
ROM_MEM[9141 ] = 8'h1B;
ROM_MEM[9142 ] = 8'h80;
ROM_MEM[9143 ] = 8'h00;
ROM_MEM[9144 ] = 8'h00;
ROM_MEM[9145 ] = 8'h80;
ROM_MEM[9146 ] = 8'h60;
ROM_MEM[9147 ] = 8'h87;
ROM_MEM[9148 ] = 8'h01;
ROM_MEM[9149 ] = 8'h82;
ROM_MEM[9150 ] = 8'h05;
ROM_MEM[9151 ] = 8'h83;
ROM_MEM[9152 ] = 8'h01;
ROM_MEM[9153 ] = 8'h8E;
ROM_MEM[9154 ] = 8'h02;
ROM_MEM[9155 ] = 8'h44;
ROM_MEM[9156 ] = 8'h16;
ROM_MEM[9157 ] = 8'h44;
ROM_MEM[9158 ] = 8'h16;
ROM_MEM[9159 ] = 8'h44;
ROM_MEM[9160 ] = 8'h14;
ROM_MEM[9161 ] = 8'h44;
ROM_MEM[9162 ] = 8'h17;
ROM_MEM[9163 ] = 8'h44;
ROM_MEM[9164 ] = 8'h16;
ROM_MEM[9165 ] = 8'h44;
ROM_MEM[9166 ] = 8'h14;
ROM_MEM[9167 ] = 8'h45;
ROM_MEM[9168 ] = 8'h16;
ROM_MEM[9169 ] = 8'h45;
ROM_MEM[9170 ] = 8'h16;
ROM_MEM[9171 ] = 8'h45;
ROM_MEM[9172 ] = 8'h14;
ROM_MEM[9173 ] = 8'h47;
ROM_MEM[9174 ] = 8'h16;
ROM_MEM[9175 ] = 8'h47;
ROM_MEM[9176 ] = 8'h16;
ROM_MEM[9177 ] = 8'h47;
ROM_MEM[9178 ] = 8'h14;
ROM_MEM[9179 ] = 8'h85;
ROM_MEM[9180 ] = 8'hF4;
ROM_MEM[9181 ] = 8'h8F;
ROM_MEM[9182 ] = 8'h00;
ROM_MEM[9183 ] = 8'h84;
ROM_MEM[9184 ] = 8'h00;
ROM_MEM[9185 ] = 8'h82;
ROM_MEM[9186 ] = 8'h07;
ROM_MEM[9187 ] = 8'h87;
ROM_MEM[9188 ] = 8'h03;
ROM_MEM[9189 ] = 8'h00;
ROM_MEM[9190 ] = 8'h80;
ROM_MEM[9191 ] = 8'h00;
ROM_MEM[9192 ] = 8'h80;
ROM_MEM[9193 ] = 8'h00;
ROM_MEM[9194 ] = 8'h80;
ROM_MEM[9195 ] = 8'h00;
ROM_MEM[9196 ] = 8'h20;
ROM_MEM[9197 ] = 8'h3F;
ROM_MEM[9198 ] = 8'h20;
ROM_MEM[9199 ] = 8'h44;
ROM_MEM[9200 ] = 8'h20;
ROM_MEM[9201 ] = 8'h49;
ROM_MEM[9202 ] = 8'h20;
ROM_MEM[9203 ] = 8'h47;
ROM_MEM[9204 ] = 8'hC0;
ROM_MEM[9205 ] = 8'h00;
ROM_MEM[9206 ] = 8'h20;
ROM_MEM[9207 ] = 8'h47;
ROM_MEM[9208 ] = 8'h20;
ROM_MEM[9209 ] = 8'h49;
ROM_MEM[9210 ] = 8'h60;
ROM_MEM[9211 ] = 8'h49;
ROM_MEM[9212 ] = 8'h20;
ROM_MEM[9213 ] = 8'h49;
ROM_MEM[9214 ] = 8'h60;
ROM_MEM[9215 ] = 8'h49;
ROM_MEM[9216 ] = 8'h20;
ROM_MEM[9217 ] = 8'h83;
ROM_MEM[9218 ] = 8'hFF;
ROM_MEM[9219 ] = 8'h87;
ROM_MEM[9220 ] = 8'h01;
ROM_MEM[9221 ] = 8'h46;
ROM_MEM[9222 ] = 8'h16;
ROM_MEM[9223 ] = 8'h46;
ROM_MEM[9224 ] = 8'h16;
ROM_MEM[9225 ] = 8'h46;
ROM_MEM[9226 ] = 8'h14;
ROM_MEM[9227 ] = 8'h46;
ROM_MEM[9228 ] = 8'h17;
ROM_MEM[9229 ] = 8'h46;
ROM_MEM[9230 ] = 8'h16;
ROM_MEM[9231 ] = 8'h46;
ROM_MEM[9232 ] = 8'h14;
ROM_MEM[9233 ] = 8'h46;
ROM_MEM[9234 ] = 8'h16;
ROM_MEM[9235 ] = 8'h00;
ROM_MEM[9236 ] = 8'h16;
ROM_MEM[9237 ] = 8'h00;
ROM_MEM[9238 ] = 8'h14;
ROM_MEM[9239 ] = 8'h00;
ROM_MEM[9240 ] = 8'h40;
ROM_MEM[9241 ] = 8'h82;
ROM_MEM[9242 ] = 8'h07;
ROM_MEM[9243 ] = 8'h87;
ROM_MEM[9244 ] = 8'h03;
ROM_MEM[9245 ] = 8'h00;
ROM_MEM[9246 ] = 8'h20;
ROM_MEM[9247 ] = 8'h44;
ROM_MEM[9248 ] = 8'h60;
ROM_MEM[9249 ] = 8'h45;
ROM_MEM[9250 ] = 8'h40;
ROM_MEM[9251 ] = 8'h47;
ROM_MEM[9252 ] = 8'h20;
ROM_MEM[9253 ] = 8'h00;
ROM_MEM[9254 ] = 8'h00;
ROM_MEM[9255 ] = 8'h80;
ROM_MEM[9256 ] = 8'h60;
ROM_MEM[9257 ] = 8'h87;
ROM_MEM[9258 ] = 8'h01;
ROM_MEM[9259 ] = 8'h82;
ROM_MEM[9260 ] = 8'h05;
ROM_MEM[9261 ] = 8'h83;
ROM_MEM[9262 ] = 8'h01;
ROM_MEM[9263 ] = 8'h8E;
ROM_MEM[9264 ] = 8'h02;
ROM_MEM[9265 ] = 8'h41;
ROM_MEM[9266 ] = 8'h16;
ROM_MEM[9267 ] = 8'h41;
ROM_MEM[9268 ] = 8'h16;
ROM_MEM[9269 ] = 8'h41;
ROM_MEM[9270 ] = 8'h14;
ROM_MEM[9271 ] = 8'h41;
ROM_MEM[9272 ] = 8'h17;
ROM_MEM[9273 ] = 8'h41;
ROM_MEM[9274 ] = 8'h16;
ROM_MEM[9275 ] = 8'h41;
ROM_MEM[9276 ] = 8'h14;
ROM_MEM[9277 ] = 8'h42;
ROM_MEM[9278 ] = 8'h16;
ROM_MEM[9279 ] = 8'h42;
ROM_MEM[9280 ] = 8'h16;
ROM_MEM[9281 ] = 8'h42;
ROM_MEM[9282 ] = 8'h14;
ROM_MEM[9283 ] = 8'h44;
ROM_MEM[9284 ] = 8'h16;
ROM_MEM[9285 ] = 8'h44;
ROM_MEM[9286 ] = 8'h16;
ROM_MEM[9287 ] = 8'h44;
ROM_MEM[9288 ] = 8'h14;
ROM_MEM[9289 ] = 8'h85;
ROM_MEM[9290 ] = 8'hF4;
ROM_MEM[9291 ] = 8'h8F;
ROM_MEM[9292 ] = 8'h00;
ROM_MEM[9293 ] = 8'h84;
ROM_MEM[9294 ] = 8'h00;
ROM_MEM[9295 ] = 8'h82;
ROM_MEM[9296 ] = 8'h07;
ROM_MEM[9297 ] = 8'h87;
ROM_MEM[9298 ] = 8'h03;
ROM_MEM[9299 ] = 8'h00;
ROM_MEM[9300 ] = 8'h60;
ROM_MEM[9301 ] = 8'h36;
ROM_MEM[9302 ] = 8'h20;
ROM_MEM[9303 ] = 8'h3B;
ROM_MEM[9304 ] = 8'h60;
ROM_MEM[9305 ] = 8'h38;
ROM_MEM[9306 ] = 8'h20;
ROM_MEM[9307 ] = 8'h3F;
ROM_MEM[9308 ] = 8'h60;
ROM_MEM[9309 ] = 8'h38;
ROM_MEM[9310 ] = 8'h20;
ROM_MEM[9311 ] = 8'h3D;
ROM_MEM[9312 ] = 8'h20;
ROM_MEM[9313 ] = 8'h42;
ROM_MEM[9314 ] = 8'h60;
ROM_MEM[9315 ] = 8'h00;
ROM_MEM[9316 ] = 8'h20;
ROM_MEM[9317 ] = 8'h3D;
ROM_MEM[9318 ] = 8'h20;
ROM_MEM[9319 ] = 8'h42;
ROM_MEM[9320 ] = 8'h20;
ROM_MEM[9321 ] = 8'h86;
ROM_MEM[9322 ] = 8'h01;
ROM_MEM[9323 ] = 8'h47;
ROM_MEM[9324 ] = 8'h20;
ROM_MEM[9325 ] = 8'h86;
ROM_MEM[9326 ] = 8'h00;
ROM_MEM[9327 ] = 8'h00;
ROM_MEM[9328 ] = 8'h20;
ROM_MEM[9329 ] = 8'h36;
ROM_MEM[9330 ] = 8'h20;
ROM_MEM[9331 ] = 8'h3B;
ROM_MEM[9332 ] = 8'h20;
ROM_MEM[9333 ] = 8'h40;
ROM_MEM[9334 ] = 8'h20;
ROM_MEM[9335 ] = 8'h3D;
ROM_MEM[9336 ] = 8'h20;
ROM_MEM[9337 ] = 8'h42;
ROM_MEM[9338 ] = 8'h20;
ROM_MEM[9339 ] = 8'h86;
ROM_MEM[9340 ] = 8'h01;
ROM_MEM[9341 ] = 8'h47;
ROM_MEM[9342 ] = 8'h20;
ROM_MEM[9343 ] = 8'h49;
ROM_MEM[9344 ] = 8'h20;
ROM_MEM[9345 ] = 8'h86;
ROM_MEM[9346 ] = 8'h00;
ROM_MEM[9347 ] = 8'h00;
ROM_MEM[9348 ] = 8'h20;
ROM_MEM[9349 ] = 8'h36;
ROM_MEM[9350 ] = 8'h20;
ROM_MEM[9351 ] = 8'h3B;
ROM_MEM[9352 ] = 8'h20;
ROM_MEM[9353 ] = 8'h40;
ROM_MEM[9354 ] = 8'h20;
ROM_MEM[9355 ] = 8'h83;
ROM_MEM[9356 ] = 8'hFF;
ROM_MEM[9357 ] = 8'h87;
ROM_MEM[9358 ] = 8'h01;
ROM_MEM[9359 ] = 8'h44;
ROM_MEM[9360 ] = 8'h16;
ROM_MEM[9361 ] = 8'h44;
ROM_MEM[9362 ] = 8'h16;
ROM_MEM[9363 ] = 8'h44;
ROM_MEM[9364 ] = 8'h14;
ROM_MEM[9365 ] = 8'h44;
ROM_MEM[9366 ] = 8'h17;
ROM_MEM[9367 ] = 8'h44;
ROM_MEM[9368 ] = 8'h16;
ROM_MEM[9369 ] = 8'h44;
ROM_MEM[9370 ] = 8'h14;
ROM_MEM[9371 ] = 8'h44;
ROM_MEM[9372 ] = 8'h16;
ROM_MEM[9373 ] = 8'h00;
ROM_MEM[9374 ] = 8'h16;
ROM_MEM[9375 ] = 8'h00;
ROM_MEM[9376 ] = 8'h14;
ROM_MEM[9377 ] = 8'h00;
ROM_MEM[9378 ] = 8'h40;
ROM_MEM[9379 ] = 8'h82;
ROM_MEM[9380 ] = 8'h07;
ROM_MEM[9381 ] = 8'h87;
ROM_MEM[9382 ] = 8'h03;
ROM_MEM[9383 ] = 8'h00;
ROM_MEM[9384 ] = 8'h20;
ROM_MEM[9385 ] = 8'h41;
ROM_MEM[9386 ] = 8'h60;
ROM_MEM[9387 ] = 8'h42;
ROM_MEM[9388 ] = 8'h40;
ROM_MEM[9389 ] = 8'h43;
ROM_MEM[9390 ] = 8'h20;
ROM_MEM[9391 ] = 8'h00;
ROM_MEM[9392 ] = 8'h00;
ROM_MEM[9393 ] = 8'h80;
ROM_MEM[9394 ] = 8'h60;
ROM_MEM[9395 ] = 8'h87;
ROM_MEM[9396 ] = 8'h01;
ROM_MEM[9397 ] = 8'h82;
ROM_MEM[9398 ] = 8'h05;
ROM_MEM[9399 ] = 8'h83;
ROM_MEM[9400 ] = 8'h01;
ROM_MEM[9401 ] = 8'h8E;
ROM_MEM[9402 ] = 8'h02;
ROM_MEM[9403 ] = 8'h3D;
ROM_MEM[9404 ] = 8'h16;
ROM_MEM[9405 ] = 8'h3D;
ROM_MEM[9406 ] = 8'h16;
ROM_MEM[9407 ] = 8'h3D;
ROM_MEM[9408 ] = 8'h14;
ROM_MEM[9409 ] = 8'h3D;
ROM_MEM[9410 ] = 8'h17;
ROM_MEM[9411 ] = 8'h3D;
ROM_MEM[9412 ] = 8'h16;
ROM_MEM[9413 ] = 8'h3D;
ROM_MEM[9414 ] = 8'h14;
ROM_MEM[9415 ] = 8'h3E;
ROM_MEM[9416 ] = 8'h16;
ROM_MEM[9417 ] = 8'h3E;
ROM_MEM[9418 ] = 8'h16;
ROM_MEM[9419 ] = 8'h3E;
ROM_MEM[9420 ] = 8'h14;
ROM_MEM[9421 ] = 8'h40;
ROM_MEM[9422 ] = 8'h16;
ROM_MEM[9423 ] = 8'h40;
ROM_MEM[9424 ] = 8'h16;
ROM_MEM[9425 ] = 8'h40;
ROM_MEM[9426 ] = 8'h14;
ROM_MEM[9427 ] = 8'h85;
ROM_MEM[9428 ] = 8'hF4;
ROM_MEM[9429 ] = 8'h8F;
ROM_MEM[9430 ] = 8'h00;
ROM_MEM[9431 ] = 8'h84;
ROM_MEM[9432 ] = 8'h00;
ROM_MEM[9433 ] = 8'h82;
ROM_MEM[9434 ] = 8'h07;
ROM_MEM[9435 ] = 8'h87;
ROM_MEM[9436 ] = 8'h03;
ROM_MEM[9437 ] = 8'h00;
ROM_MEM[9438 ] = 8'h20;
ROM_MEM[9439 ] = 8'h2C;
ROM_MEM[9440 ] = 8'h20;
ROM_MEM[9441 ] = 8'h31;
ROM_MEM[9442 ] = 8'h60;
ROM_MEM[9443 ] = 8'h2F;
ROM_MEM[9444 ] = 8'h20;
ROM_MEM[9445 ] = 8'h34;
ROM_MEM[9446 ] = 8'h40;
ROM_MEM[9447 ] = 8'h00;
ROM_MEM[9448 ] = 8'h20;
ROM_MEM[9449 ] = 8'h2C;
ROM_MEM[9450 ] = 8'h20;
ROM_MEM[9451 ] = 8'h31;
ROM_MEM[9452 ] = 8'h20;
ROM_MEM[9453 ] = 8'h36;
ROM_MEM[9454 ] = 8'h20;
ROM_MEM[9455 ] = 8'h33;
ROM_MEM[9456 ] = 8'h20;
ROM_MEM[9457 ] = 8'h2E;
ROM_MEM[9458 ] = 8'h20;
ROM_MEM[9459 ] = 8'h31;
ROM_MEM[9460 ] = 8'h20;
ROM_MEM[9461 ] = 8'h2C;
ROM_MEM[9462 ] = 8'h40;
ROM_MEM[9463 ] = 8'h31;
ROM_MEM[9464 ] = 8'h20;
ROM_MEM[9465 ] = 8'h2C;
ROM_MEM[9466 ] = 8'h20;
ROM_MEM[9467 ] = 8'h27;
ROM_MEM[9468 ] = 8'h40;
ROM_MEM[9469 ] = 8'h2C;
ROM_MEM[9470 ] = 8'h20;
ROM_MEM[9471 ] = 8'h27;
ROM_MEM[9472 ] = 8'h20;
ROM_MEM[9473 ] = 8'h22;
ROM_MEM[9474 ] = 8'h20;
ROM_MEM[9475 ] = 8'h00;
ROM_MEM[9476 ] = 8'h20;
ROM_MEM[9477 ] = 8'h34;
ROM_MEM[9478 ] = 8'h20;
ROM_MEM[9479 ] = 8'h2F;
ROM_MEM[9480 ] = 8'h20;
ROM_MEM[9481 ] = 8'h2A;
ROM_MEM[9482 ] = 8'h20;
ROM_MEM[9483 ] = 8'h00;
ROM_MEM[9484 ] = 8'h20;
ROM_MEM[9485 ] = 8'h2F;
ROM_MEM[9486 ] = 8'h20;
ROM_MEM[9487 ] = 8'h2A;
ROM_MEM[9488 ] = 8'h20;
ROM_MEM[9489 ] = 8'h25;
ROM_MEM[9490 ] = 8'h20;
ROM_MEM[9491 ] = 8'h83;
ROM_MEM[9492 ] = 8'hFF;
ROM_MEM[9493 ] = 8'h87;
ROM_MEM[9494 ] = 8'h01;
ROM_MEM[9495 ] = 8'h3F;
ROM_MEM[9496 ] = 8'h16;
ROM_MEM[9497 ] = 8'h3F;
ROM_MEM[9498 ] = 8'h16;
ROM_MEM[9499 ] = 8'h3F;
ROM_MEM[9500 ] = 8'h14;
ROM_MEM[9501 ] = 8'h3F;
ROM_MEM[9502 ] = 8'h17;
ROM_MEM[9503 ] = 8'h3F;
ROM_MEM[9504 ] = 8'h16;
ROM_MEM[9505 ] = 8'h3F;
ROM_MEM[9506 ] = 8'h14;
ROM_MEM[9507 ] = 8'h3F;
ROM_MEM[9508 ] = 8'h16;
ROM_MEM[9509 ] = 8'h2E;
ROM_MEM[9510 ] = 8'h16;
ROM_MEM[9511 ] = 8'h33;
ROM_MEM[9512 ] = 8'h14;
ROM_MEM[9513 ] = 8'h38;
ROM_MEM[9514 ] = 8'h16;
ROM_MEM[9515 ] = 8'h3A;
ROM_MEM[9516 ] = 8'h16;
ROM_MEM[9517 ] = 8'h3B;
ROM_MEM[9518 ] = 8'h14;
ROM_MEM[9519 ] = 8'h82;
ROM_MEM[9520 ] = 8'h07;
ROM_MEM[9521 ] = 8'h87;
ROM_MEM[9522 ] = 8'h03;
ROM_MEM[9523 ] = 8'h00;
ROM_MEM[9524 ] = 8'h20;
ROM_MEM[9525 ] = 8'h31;
ROM_MEM[9526 ] = 8'h10;
ROM_MEM[9527 ] = 8'h35;
ROM_MEM[9528 ] = 8'h10;
ROM_MEM[9529 ] = 8'h39;
ROM_MEM[9530 ] = 8'h16;
ROM_MEM[9531 ] = 8'h3D;
ROM_MEM[9532 ] = 8'h16;
ROM_MEM[9533 ] = 8'h86;
ROM_MEM[9534 ] = 8'h01;
ROM_MEM[9535 ] = 8'h41;
ROM_MEM[9536 ] = 8'h14;
ROM_MEM[9537 ] = 8'h42;
ROM_MEM[9538 ] = 8'h16;
ROM_MEM[9539 ] = 8'h44;
ROM_MEM[9540 ] = 8'h16;
ROM_MEM[9541 ] = 8'h45;
ROM_MEM[9542 ] = 8'h14;
ROM_MEM[9543 ] = 8'h86;
ROM_MEM[9544 ] = 8'h00;
ROM_MEM[9545 ] = 8'h40;
ROM_MEM[9546 ] = 8'h20;
ROM_MEM[9547 ] = 8'h00;
ROM_MEM[9548 ] = 8'h00;
ROM_MEM[9549 ] = 8'h80;
ROM_MEM[9550 ] = 8'h60;
ROM_MEM[9551 ] = 8'h87;
ROM_MEM[9552 ] = 8'h01;
ROM_MEM[9553 ] = 8'h2D;
ROM_MEM[9554 ] = 8'h16;
ROM_MEM[9555 ] = 8'h2D;
ROM_MEM[9556 ] = 8'h16;
ROM_MEM[9557 ] = 8'h2D;
ROM_MEM[9558 ] = 8'h14;
ROM_MEM[9559 ] = 8'h2D;
ROM_MEM[9560 ] = 8'h17;
ROM_MEM[9561 ] = 8'h2D;
ROM_MEM[9562 ] = 8'h16;
ROM_MEM[9563 ] = 8'h2D;
ROM_MEM[9564 ] = 8'h14;
ROM_MEM[9565 ] = 8'h2C;
ROM_MEM[9566 ] = 8'h16;
ROM_MEM[9567 ] = 8'h2C;
ROM_MEM[9568 ] = 8'h16;
ROM_MEM[9569 ] = 8'h2C;
ROM_MEM[9570 ] = 8'h14;
ROM_MEM[9571 ] = 8'h2A;
ROM_MEM[9572 ] = 8'h16;
ROM_MEM[9573 ] = 8'h2A;
ROM_MEM[9574 ] = 8'h16;
ROM_MEM[9575 ] = 8'h2A;
ROM_MEM[9576 ] = 8'h14;
ROM_MEM[9577 ] = 8'h21;
ROM_MEM[9578 ] = 8'h16;
ROM_MEM[9579 ] = 8'h21;
ROM_MEM[9580 ] = 8'h16;
ROM_MEM[9581 ] = 8'h21;
ROM_MEM[9582 ] = 8'h14;
ROM_MEM[9583 ] = 8'h21;
ROM_MEM[9584 ] = 8'h17;
ROM_MEM[9585 ] = 8'h21;
ROM_MEM[9586 ] = 8'h16;
ROM_MEM[9587 ] = 8'h21;
ROM_MEM[9588 ] = 8'h14;
ROM_MEM[9589 ] = 8'h20;
ROM_MEM[9590 ] = 8'h16;
ROM_MEM[9591 ] = 8'h20;
ROM_MEM[9592 ] = 8'h16;
ROM_MEM[9593 ] = 8'h1E;
ROM_MEM[9594 ] = 8'h14;
ROM_MEM[9595 ] = 8'h1D;
ROM_MEM[9596 ] = 8'h16;
ROM_MEM[9597 ] = 8'h1D;
ROM_MEM[9598 ] = 8'h16;
ROM_MEM[9599 ] = 8'h1D;
ROM_MEM[9600 ] = 8'h14;
ROM_MEM[9601 ] = 8'h87;
ROM_MEM[9602 ] = 8'h03;
ROM_MEM[9603 ] = 8'h25;
ROM_MEM[9604 ] = 8'h40;
ROM_MEM[9605 ] = 8'h00;
ROM_MEM[9606 ] = 8'h40;
ROM_MEM[9607 ] = 8'h00;
ROM_MEM[9608 ] = 8'h80;
ROM_MEM[9609 ] = 8'h00;
ROM_MEM[9610 ] = 8'h80;
ROM_MEM[9611 ] = 8'h00;
ROM_MEM[9612 ] = 8'h80;
ROM_MEM[9613 ] = 8'h00;
ROM_MEM[9614 ] = 8'h20;
ROM_MEM[9615 ] = 8'h86;
ROM_MEM[9616 ] = 8'h01;
ROM_MEM[9617 ] = 8'h31;
ROM_MEM[9618 ] = 8'h60;
ROM_MEM[9619 ] = 8'h86;
ROM_MEM[9620 ] = 8'h00;
ROM_MEM[9621 ] = 8'h2F;
ROM_MEM[9622 ] = 8'h20;
ROM_MEM[9623 ] = 8'h34;
ROM_MEM[9624 ] = 8'h20;
ROM_MEM[9625 ] = 8'h31;
ROM_MEM[9626 ] = 8'h20;
ROM_MEM[9627 ] = 8'h36;
ROM_MEM[9628 ] = 8'h20;
ROM_MEM[9629 ] = 8'h47;
ROM_MEM[9630 ] = 8'h60;
ROM_MEM[9631 ] = 8'h47;
ROM_MEM[9632 ] = 8'h20;
ROM_MEM[9633 ] = 8'h47;
ROM_MEM[9634 ] = 8'h60;
ROM_MEM[9635 ] = 8'h47;
ROM_MEM[9636 ] = 8'h20;
ROM_MEM[9637 ] = 8'h87;
ROM_MEM[9638 ] = 8'h01;
ROM_MEM[9639 ] = 8'h2E;
ROM_MEM[9640 ] = 8'h16;
ROM_MEM[9641 ] = 8'h2E;
ROM_MEM[9642 ] = 8'h16;
ROM_MEM[9643 ] = 8'h2E;
ROM_MEM[9644 ] = 8'h14;
ROM_MEM[9645 ] = 8'h2E;
ROM_MEM[9646 ] = 8'h17;
ROM_MEM[9647 ] = 8'h2E;
ROM_MEM[9648 ] = 8'h16;
ROM_MEM[9649 ] = 8'h2E;
ROM_MEM[9650 ] = 8'h14;
ROM_MEM[9651 ] = 8'h2E;
ROM_MEM[9652 ] = 8'h16;
ROM_MEM[9653 ] = 8'h27;
ROM_MEM[9654 ] = 8'h16;
ROM_MEM[9655 ] = 8'h22;
ROM_MEM[9656 ] = 8'h14;
ROM_MEM[9657 ] = 8'h1D;
ROM_MEM[9658 ] = 8'h16;
ROM_MEM[9659 ] = 8'h1B;
ROM_MEM[9660 ] = 8'h16;
ROM_MEM[9661 ] = 8'h1A;
ROM_MEM[9662 ] = 8'h14;
ROM_MEM[9663 ] = 8'h87;
ROM_MEM[9664 ] = 8'h03;
ROM_MEM[9665 ] = 8'h00;
ROM_MEM[9666 ] = 8'h20;
ROM_MEM[9667 ] = 8'h2D;
ROM_MEM[9668 ] = 8'h60;
ROM_MEM[9669 ] = 8'h2C;
ROM_MEM[9670 ] = 8'h40;
ROM_MEM[9671 ] = 8'h25;
ROM_MEM[9672 ] = 8'h20;
ROM_MEM[9673 ] = 8'h00;
ROM_MEM[9674 ] = 8'h00;
ROM_MEM[9675 ] = 8'h80;
ROM_MEM[9676 ] = 8'h80;
ROM_MEM[9677 ] = 8'h87;
ROM_MEM[9678 ] = 8'h03;
ROM_MEM[9679 ] = 8'h36;
ROM_MEM[9680 ] = 8'h2A;
ROM_MEM[9681 ] = 8'h36;
ROM_MEM[9682 ] = 8'h2A;
ROM_MEM[9683 ] = 8'h36;
ROM_MEM[9684 ] = 8'h2C;
ROM_MEM[9685 ] = 8'h3B;
ROM_MEM[9686 ] = 8'h80;
ROM_MEM[9687 ] = 8'h3B;
ROM_MEM[9688 ] = 8'h81;
ROM_MEM[9689 ] = 8'h42;
ROM_MEM[9690 ] = 8'hC0;
ROM_MEM[9691 ] = 8'h42;
ROM_MEM[9692 ] = 8'h21;
ROM_MEM[9693 ] = 8'h00;
ROM_MEM[9694 ] = 8'h20;
ROM_MEM[9695 ] = 8'h8E;
ROM_MEM[9696 ] = 8'h02;
ROM_MEM[9697 ] = 8'h40;
ROM_MEM[9698 ] = 8'h16;
ROM_MEM[9699 ] = 8'h3F;
ROM_MEM[9700 ] = 8'h16;
ROM_MEM[9701 ] = 8'h3D;
ROM_MEM[9702 ] = 8'h14;
ROM_MEM[9703 ] = 8'h47;
ROM_MEM[9704 ] = 8'hC0;
ROM_MEM[9705 ] = 8'h42;
ROM_MEM[9706 ] = 8'hC0;
ROM_MEM[9707 ] = 8'h42;
ROM_MEM[9708 ] = 8'h21;
ROM_MEM[9709 ] = 8'h00;
ROM_MEM[9710 ] = 8'h20;
ROM_MEM[9711 ] = 8'h8F;
ROM_MEM[9712 ] = 8'h00;
ROM_MEM[9713 ] = 8'h40;
ROM_MEM[9714 ] = 8'h16;
ROM_MEM[9715 ] = 8'h3F;
ROM_MEM[9716 ] = 8'h16;
ROM_MEM[9717 ] = 8'h40;
ROM_MEM[9718 ] = 8'h14;
ROM_MEM[9719 ] = 8'h3D;
ROM_MEM[9720 ] = 8'hC0;
ROM_MEM[9721 ] = 8'h3D;
ROM_MEM[9722 ] = 8'hC1;
ROM_MEM[9723 ] = 8'h00;
ROM_MEM[9724 ] = 8'h00;
ROM_MEM[9725 ] = 8'h80;
ROM_MEM[9726 ] = 8'h80;
ROM_MEM[9727 ] = 8'h87;
ROM_MEM[9728 ] = 8'h03;
ROM_MEM[9729 ] = 8'h2A;
ROM_MEM[9730 ] = 8'h2A;
ROM_MEM[9731 ] = 8'h2A;
ROM_MEM[9732 ] = 8'h2A;
ROM_MEM[9733 ] = 8'h2A;
ROM_MEM[9734 ] = 8'h2C;
ROM_MEM[9735 ] = 8'h33;
ROM_MEM[9736 ] = 8'h80;
ROM_MEM[9737 ] = 8'h33;
ROM_MEM[9738 ] = 8'h81;
ROM_MEM[9739 ] = 8'h3B;
ROM_MEM[9740 ] = 8'hC0;
ROM_MEM[9741 ] = 8'h3B;
ROM_MEM[9742 ] = 8'h21;
ROM_MEM[9743 ] = 8'h00;
ROM_MEM[9744 ] = 8'h20;
ROM_MEM[9745 ] = 8'h8E;
ROM_MEM[9746 ] = 8'h02;
ROM_MEM[9747 ] = 8'h38;
ROM_MEM[9748 ] = 8'h40;
ROM_MEM[9749 ] = 8'h3F;
ROM_MEM[9750 ] = 8'hC0;
ROM_MEM[9751 ] = 8'h3B;
ROM_MEM[9752 ] = 8'hC0;
ROM_MEM[9753 ] = 8'h3B;
ROM_MEM[9754 ] = 8'h21;
ROM_MEM[9755 ] = 8'h00;
ROM_MEM[9756 ] = 8'h20;
ROM_MEM[9757 ] = 8'h8F;
ROM_MEM[9758 ] = 8'h00;
ROM_MEM[9759 ] = 8'h3D;
ROM_MEM[9760 ] = 8'h16;
ROM_MEM[9761 ] = 8'h3C;
ROM_MEM[9762 ] = 8'h16;
ROM_MEM[9763 ] = 8'h3D;
ROM_MEM[9764 ] = 8'h14;
ROM_MEM[9765 ] = 8'h39;
ROM_MEM[9766 ] = 8'hC0;
ROM_MEM[9767 ] = 8'h3A;
ROM_MEM[9768 ] = 8'hC0;
ROM_MEM[9769 ] = 8'h00;
ROM_MEM[9770 ] = 8'h00;
ROM_MEM[9771 ] = 8'h80;
ROM_MEM[9772 ] = 8'h80;
ROM_MEM[9773 ] = 8'h87;
ROM_MEM[9774 ] = 8'h03;
ROM_MEM[9775 ] = 8'h00;
ROM_MEM[9776 ] = 8'h80;
ROM_MEM[9777 ] = 8'h8E;
ROM_MEM[9778 ] = 8'h0E;
ROM_MEM[9779 ] = 8'h20;
ROM_MEM[9780 ] = 8'h40;
ROM_MEM[9781 ] = 8'h20;
ROM_MEM[9782 ] = 8'h40;
ROM_MEM[9783 ] = 8'h8F;
ROM_MEM[9784 ] = 8'h00;
ROM_MEM[9785 ] = 8'h2A;
ROM_MEM[9786 ] = 8'hC0;
ROM_MEM[9787 ] = 8'h00;
ROM_MEM[9788 ] = 8'h00;
ROM_MEM[9789 ] = 8'h80;
ROM_MEM[9790 ] = 8'h80;
ROM_MEM[9791 ] = 8'h87;
ROM_MEM[9792 ] = 8'h04;
ROM_MEM[9793 ] = 8'h82;
ROM_MEM[9794 ] = 8'h0A;
ROM_MEM[9795 ] = 8'h1E;
ROM_MEM[9796 ] = 8'h2A;
ROM_MEM[9797 ] = 8'h1E;
ROM_MEM[9798 ] = 8'h2A;
ROM_MEM[9799 ] = 8'h1E;
ROM_MEM[9800 ] = 8'h2C;
ROM_MEM[9801 ] = 8'h00;
ROM_MEM[9802 ] = 8'h80;
ROM_MEM[9803 ] = 8'h25;
ROM_MEM[9804 ] = 8'h80;
ROM_MEM[9805 ] = 8'h25;
ROM_MEM[9806 ] = 8'h81;
ROM_MEM[9807 ] = 8'h27;
ROM_MEM[9808 ] = 8'h80;
ROM_MEM[9809 ] = 8'h27;
ROM_MEM[9810 ] = 8'h81;
ROM_MEM[9811 ] = 8'h28;
ROM_MEM[9812 ] = 8'h80;
ROM_MEM[9813 ] = 8'h28;
ROM_MEM[9814 ] = 8'h81;
ROM_MEM[9815 ] = 8'h2A;
ROM_MEM[9816 ] = 8'h80;
ROM_MEM[9817 ] = 8'h2A;
ROM_MEM[9818 ] = 8'h81;
ROM_MEM[9819 ] = 8'h2C;
ROM_MEM[9820 ] = 8'h80;
ROM_MEM[9821 ] = 8'h2C;
ROM_MEM[9822 ] = 8'h81;
ROM_MEM[9823 ] = 8'h2E;
ROM_MEM[9824 ] = 8'h40;
ROM_MEM[9825 ] = 8'h2F;
ROM_MEM[9826 ] = 8'h40;
ROM_MEM[9827 ] = 8'h2D;
ROM_MEM[9828 ] = 8'h80;
ROM_MEM[9829 ] = 8'h2D;
ROM_MEM[9830 ] = 8'h81;
ROM_MEM[9831 ] = 8'h1E;
ROM_MEM[9832 ] = 8'hC0;
ROM_MEM[9833 ] = 8'h00;
ROM_MEM[9834 ] = 8'h00;
ROM_MEM[9835 ] = 8'h80;
ROM_MEM[9836 ] = 8'h50;
ROM_MEM[9837 ] = 8'h87;
ROM_MEM[9838 ] = 8'h02;
ROM_MEM[9839 ] = 8'h82;
ROM_MEM[9840 ] = 8'h05;
ROM_MEM[9841 ] = 8'h44;
ROM_MEM[9842 ] = 8'h16;
ROM_MEM[9843 ] = 8'h43;
ROM_MEM[9844 ] = 8'h16;
ROM_MEM[9845 ] = 8'h41;
ROM_MEM[9846 ] = 8'h14;
ROM_MEM[9847 ] = 8'h46;
ROM_MEM[9848 ] = 8'h40;
ROM_MEM[9849 ] = 8'h46;
ROM_MEM[9850 ] = 8'h17;
ROM_MEM[9851 ] = 8'h44;
ROM_MEM[9852 ] = 8'h16;
ROM_MEM[9853 ] = 8'h43;
ROM_MEM[9854 ] = 8'h14;
ROM_MEM[9855 ] = 8'h48;
ROM_MEM[9856 ] = 8'h40;
ROM_MEM[9857 ] = 8'h48;
ROM_MEM[9858 ] = 8'h17;
ROM_MEM[9859 ] = 8'h46;
ROM_MEM[9860 ] = 8'h16;
ROM_MEM[9861 ] = 8'h44;
ROM_MEM[9862 ] = 8'h14;
ROM_MEM[9863 ] = 8'h49;
ROM_MEM[9864 ] = 8'h16;
ROM_MEM[9865 ] = 8'h48;
ROM_MEM[9866 ] = 8'h16;
ROM_MEM[9867 ] = 8'h46;
ROM_MEM[9868 ] = 8'h14;
ROM_MEM[9869 ] = 8'h4D;
ROM_MEM[9870 ] = 8'h16;
ROM_MEM[9871 ] = 8'h4B;
ROM_MEM[9872 ] = 8'h16;
ROM_MEM[9873 ] = 8'h49;
ROM_MEM[9874 ] = 8'h14;
ROM_MEM[9875 ] = 8'h4F;
ROM_MEM[9876 ] = 8'h16;
ROM_MEM[9877 ] = 8'h4D;
ROM_MEM[9878 ] = 8'h16;
ROM_MEM[9879 ] = 8'h4B;
ROM_MEM[9880 ] = 8'h14;
ROM_MEM[9881 ] = 8'h82;
ROM_MEM[9882 ] = 8'h03;
ROM_MEM[9883 ] = 8'h50;
ROM_MEM[9884 ] = 8'h80;
ROM_MEM[9885 ] = 8'h50;
ROM_MEM[9886 ] = 8'h81;
ROM_MEM[9887 ] = 8'h82;
ROM_MEM[9888 ] = 8'h07;
ROM_MEM[9889 ] = 8'h87;
ROM_MEM[9890 ] = 8'h03;
ROM_MEM[9891 ] = 8'h3F;
ROM_MEM[9892 ] = 8'h20;
ROM_MEM[9893 ] = 8'h00;
ROM_MEM[9894 ] = 8'h20;
ROM_MEM[9895 ] = 8'h3F;
ROM_MEM[9896 ] = 8'h16;
ROM_MEM[9897 ] = 8'h3F;
ROM_MEM[9898 ] = 8'h16;
ROM_MEM[9899 ] = 8'h3F;
ROM_MEM[9900 ] = 8'h14;
ROM_MEM[9901 ] = 8'h3F;
ROM_MEM[9902 ] = 8'h40;
ROM_MEM[9903 ] = 8'h00;
ROM_MEM[9904 ] = 8'h00;
ROM_MEM[9905 ] = 8'h80;
ROM_MEM[9906 ] = 8'h50;
ROM_MEM[9907 ] = 8'h87;
ROM_MEM[9908 ] = 8'h03;
ROM_MEM[9909 ] = 8'h00;
ROM_MEM[9910 ] = 8'h40;
ROM_MEM[9911 ] = 8'h41;
ROM_MEM[9912 ] = 8'h80;
ROM_MEM[9913 ] = 8'h41;
ROM_MEM[9914 ] = 8'h80;
ROM_MEM[9915 ] = 8'h41;
ROM_MEM[9916 ] = 8'h80;
ROM_MEM[9917 ] = 8'h41;
ROM_MEM[9918 ] = 8'h40;
ROM_MEM[9919 ] = 8'h82;
ROM_MEM[9920 ] = 8'h09;
ROM_MEM[9921 ] = 8'h44;
ROM_MEM[9922 ] = 8'h20;
ROM_MEM[9923 ] = 8'h42;
ROM_MEM[9924 ] = 8'h20;
ROM_MEM[9925 ] = 8'h40;
ROM_MEM[9926 ] = 8'h16;
ROM_MEM[9927 ] = 8'h40;
ROM_MEM[9928 ] = 8'h17;
ROM_MEM[9929 ] = 8'h3F;
ROM_MEM[9930 ] = 8'h14;
ROM_MEM[9931 ] = 8'h3D;
ROM_MEM[9932 ] = 8'h20;
ROM_MEM[9933 ] = 8'h3B;
ROM_MEM[9934 ] = 8'h20;
ROM_MEM[9935 ] = 8'h3A;
ROM_MEM[9936 ] = 8'h16;
ROM_MEM[9937 ] = 8'h3A;
ROM_MEM[9938 ] = 8'h17;
ROM_MEM[9939 ] = 8'h38;
ROM_MEM[9940 ] = 8'h14;
ROM_MEM[9941 ] = 8'h82;
ROM_MEM[9942 ] = 8'h07;
ROM_MEM[9943 ] = 8'h38;
ROM_MEM[9944 ] = 8'h80;
ROM_MEM[9945 ] = 8'h37;
ROM_MEM[9946 ] = 8'h40;
ROM_MEM[9947 ] = 8'h00;
ROM_MEM[9948 ] = 8'h00;
ROM_MEM[9949 ] = 8'h80;
ROM_MEM[9950 ] = 8'h50;
ROM_MEM[9951 ] = 8'h87;
ROM_MEM[9952 ] = 8'h03;
ROM_MEM[9953 ] = 8'h00;
ROM_MEM[9954 ] = 8'h40;
ROM_MEM[9955 ] = 8'h3C;
ROM_MEM[9956 ] = 8'h80;
ROM_MEM[9957 ] = 8'h3C;
ROM_MEM[9958 ] = 8'h80;
ROM_MEM[9959 ] = 8'h3C;
ROM_MEM[9960 ] = 8'h80;
ROM_MEM[9961 ] = 8'h3C;
ROM_MEM[9962 ] = 8'h40;
ROM_MEM[9963 ] = 8'h82;
ROM_MEM[9964 ] = 8'h09;
ROM_MEM[9965 ] = 8'h40;
ROM_MEM[9966 ] = 8'h20;
ROM_MEM[9967 ] = 8'h3F;
ROM_MEM[9968 ] = 8'h20;
ROM_MEM[9969 ] = 8'h3D;
ROM_MEM[9970 ] = 8'h16;
ROM_MEM[9971 ] = 8'h3D;
ROM_MEM[9972 ] = 8'h17;
ROM_MEM[9973 ] = 8'h3B;
ROM_MEM[9974 ] = 8'h14;
ROM_MEM[9975 ] = 8'h3A;
ROM_MEM[9976 ] = 8'h20;
ROM_MEM[9977 ] = 8'h38;
ROM_MEM[9978 ] = 8'h20;
ROM_MEM[9979 ] = 8'h36;
ROM_MEM[9980 ] = 8'h16;
ROM_MEM[9981 ] = 8'h36;
ROM_MEM[9982 ] = 8'h17;
ROM_MEM[9983 ] = 8'h34;
ROM_MEM[9984 ] = 8'h14;
ROM_MEM[9985 ] = 8'h82;
ROM_MEM[9986 ] = 8'h07;
ROM_MEM[9987 ] = 8'h33;
ROM_MEM[9988 ] = 8'hC0;
ROM_MEM[9989 ] = 8'h00;
ROM_MEM[9990 ] = 8'h00;
ROM_MEM[9991 ] = 8'h80;
ROM_MEM[9992 ] = 8'h50;
ROM_MEM[9993 ] = 8'h87;
ROM_MEM[9994 ] = 8'h02;
ROM_MEM[9995 ] = 8'h00;
ROM_MEM[9996 ] = 8'h40;
ROM_MEM[9997 ] = 8'h29;
ROM_MEM[9998 ] = 8'h40;
ROM_MEM[9999 ] = 8'h2B;
ROM_MEM[10000] = 8'h40;
ROM_MEM[10001] = 8'h2C;
ROM_MEM[10002] = 8'h40;
ROM_MEM[10003] = 8'h25;
ROM_MEM[10004] = 8'h40;
ROM_MEM[10005] = 8'h2E;
ROM_MEM[10006] = 8'h40;
ROM_MEM[10007] = 8'h31;
ROM_MEM[10008] = 8'h40;
ROM_MEM[10009] = 8'h27;
ROM_MEM[10010] = 8'h40;
ROM_MEM[10011] = 8'h85;
ROM_MEM[10012] = 8'h0C;
ROM_MEM[10013] = 8'h87;
ROM_MEM[10014] = 8'h03;
ROM_MEM[10015] = 8'h16;
ROM_MEM[10016] = 8'h20;
ROM_MEM[10017] = 8'h18;
ROM_MEM[10018] = 8'h20;
ROM_MEM[10019] = 8'h19;
ROM_MEM[10020] = 8'h16;
ROM_MEM[10021] = 8'h19;
ROM_MEM[10022] = 8'h17;
ROM_MEM[10023] = 8'h1B;
ROM_MEM[10024] = 8'h14;
ROM_MEM[10025] = 8'h1C;
ROM_MEM[10026] = 8'h20;
ROM_MEM[10027] = 8'h1E;
ROM_MEM[10028] = 8'h20;
ROM_MEM[10029] = 8'h20;
ROM_MEM[10030] = 8'h16;
ROM_MEM[10031] = 8'h20;
ROM_MEM[10032] = 8'h17;
ROM_MEM[10033] = 8'h22;
ROM_MEM[10034] = 8'h14;
ROM_MEM[10035] = 8'h84;
ROM_MEM[10036] = 8'h00;
ROM_MEM[10037] = 8'h27;
ROM_MEM[10038] = 8'h20;
ROM_MEM[10039] = 8'h00;
ROM_MEM[10040] = 8'h20;
ROM_MEM[10041] = 8'h27;
ROM_MEM[10042] = 8'h16;
ROM_MEM[10043] = 8'h27;
ROM_MEM[10044] = 8'h16;
ROM_MEM[10045] = 8'h27;
ROM_MEM[10046] = 8'h14;
ROM_MEM[10047] = 8'h1B;
ROM_MEM[10048] = 8'h40;
ROM_MEM[10049] = 8'h00;
ROM_MEM[10050] = 8'h00;
ROM_MEM[10051] = 8'h82;
ROM_MEM[10052] = 8'h09;
ROM_MEM[10053] = 8'h80;
ROM_MEM[10054] = 8'h48;
ROM_MEM[10055] = 8'h87;
ROM_MEM[10056] = 8'h03;
ROM_MEM[10057] = 8'h38;
ROM_MEM[10058] = 8'h40;
ROM_MEM[10059] = 8'h38;
ROM_MEM[10060] = 8'h40;
ROM_MEM[10061] = 8'h8E;
ROM_MEM[10062] = 8'h02;
ROM_MEM[10063] = 8'h38;
ROM_MEM[10064] = 8'h40;
ROM_MEM[10065] = 8'h34;
ROM_MEM[10066] = 8'h30;
ROM_MEM[10067] = 8'h3B;
ROM_MEM[10068] = 8'h10;
ROM_MEM[10069] = 8'h8F;
ROM_MEM[10070] = 8'h00;
ROM_MEM[10071] = 8'h38;
ROM_MEM[10072] = 8'h80;
ROM_MEM[10073] = 8'h3F;
ROM_MEM[10074] = 8'h40;
ROM_MEM[10075] = 8'h3F;
ROM_MEM[10076] = 8'h40;
ROM_MEM[10077] = 8'h3F;
ROM_MEM[10078] = 8'h40;
ROM_MEM[10079] = 8'h40;
ROM_MEM[10080] = 8'h30;
ROM_MEM[10081] = 8'h3B;
ROM_MEM[10082] = 8'h10;
ROM_MEM[10083] = 8'h37;
ROM_MEM[10084] = 8'h40;
ROM_MEM[10085] = 8'h34;
ROM_MEM[10086] = 8'h30;
ROM_MEM[10087] = 8'h3B;
ROM_MEM[10088] = 8'h10;
ROM_MEM[10089] = 8'h38;
ROM_MEM[10090] = 8'h60;
ROM_MEM[10091] = 8'h83;
ROM_MEM[10092] = 8'hFF;
ROM_MEM[10093] = 8'h38;
ROM_MEM[10094] = 8'h11;
ROM_MEM[10095] = 8'h83;
ROM_MEM[10096] = 8'hFF;
ROM_MEM[10097] = 8'h38;
ROM_MEM[10098] = 8'h11;
ROM_MEM[10099] = 8'h00;
ROM_MEM[10100] = 8'h00;
ROM_MEM[10101] = 8'h82;
ROM_MEM[10102] = 8'h09;
ROM_MEM[10103] = 8'h80;
ROM_MEM[10104] = 8'h48;
ROM_MEM[10105] = 8'h87;
ROM_MEM[10106] = 8'h03;
ROM_MEM[10107] = 8'h33;
ROM_MEM[10108] = 8'h40;
ROM_MEM[10109] = 8'h33;
ROM_MEM[10110] = 8'h40;
ROM_MEM[10111] = 8'h8E;
ROM_MEM[10112] = 8'h02;
ROM_MEM[10113] = 8'h33;
ROM_MEM[10114] = 8'h40;
ROM_MEM[10115] = 8'h2F;
ROM_MEM[10116] = 8'h30;
ROM_MEM[10117] = 8'h34;
ROM_MEM[10118] = 8'h10;
ROM_MEM[10119] = 8'h8F;
ROM_MEM[10120] = 8'h00;
ROM_MEM[10121] = 8'h33;
ROM_MEM[10122] = 8'h80;
ROM_MEM[10123] = 8'h33;
ROM_MEM[10124] = 8'h40;
ROM_MEM[10125] = 8'h33;
ROM_MEM[10126] = 8'h40;
ROM_MEM[10127] = 8'h33;
ROM_MEM[10128] = 8'h40;
ROM_MEM[10129] = 8'h34;
ROM_MEM[10130] = 8'h30;
ROM_MEM[10131] = 8'h2F;
ROM_MEM[10132] = 8'h10;
ROM_MEM[10133] = 8'h34;
ROM_MEM[10134] = 8'h40;
ROM_MEM[10135] = 8'h2F;
ROM_MEM[10136] = 8'h30;
ROM_MEM[10137] = 8'h34;
ROM_MEM[10138] = 8'h10;
ROM_MEM[10139] = 8'h33;
ROM_MEM[10140] = 8'h60;
ROM_MEM[10141] = 8'h83;
ROM_MEM[10142] = 8'hFF;
ROM_MEM[10143] = 8'h33;
ROM_MEM[10144] = 8'h11;
ROM_MEM[10145] = 8'h83;
ROM_MEM[10146] = 8'hFF;
ROM_MEM[10147] = 8'h33;
ROM_MEM[10148] = 8'h11;
ROM_MEM[10149] = 8'h00;
ROM_MEM[10150] = 8'h00;
ROM_MEM[10151] = 8'h82;
ROM_MEM[10152] = 8'h09;
ROM_MEM[10153] = 8'h80;
ROM_MEM[10154] = 8'h48;
ROM_MEM[10155] = 8'h87;
ROM_MEM[10156] = 8'h03;
ROM_MEM[10157] = 8'h2F;
ROM_MEM[10158] = 8'h40;
ROM_MEM[10159] = 8'h2F;
ROM_MEM[10160] = 8'h40;
ROM_MEM[10161] = 8'h8E;
ROM_MEM[10162] = 8'h02;
ROM_MEM[10163] = 8'h2F;
ROM_MEM[10164] = 8'h40;
ROM_MEM[10165] = 8'h2B;
ROM_MEM[10166] = 8'h40;
ROM_MEM[10167] = 8'h8F;
ROM_MEM[10168] = 8'h00;
ROM_MEM[10169] = 8'h2F;
ROM_MEM[10170] = 8'h80;
ROM_MEM[10171] = 8'h3B;
ROM_MEM[10172] = 8'h40;
ROM_MEM[10173] = 8'h3B;
ROM_MEM[10174] = 8'h40;
ROM_MEM[10175] = 8'h3B;
ROM_MEM[10176] = 8'h40;
ROM_MEM[10177] = 8'h37;
ROM_MEM[10178] = 8'h40;
ROM_MEM[10179] = 8'h2F;
ROM_MEM[10180] = 8'h40;
ROM_MEM[10181] = 8'h2B;
ROM_MEM[10182] = 8'h40;
ROM_MEM[10183] = 8'h2F;
ROM_MEM[10184] = 8'h60;
ROM_MEM[10185] = 8'h83;
ROM_MEM[10186] = 8'hFF;
ROM_MEM[10187] = 8'h2F;
ROM_MEM[10188] = 8'h11;
ROM_MEM[10189] = 8'h83;
ROM_MEM[10190] = 8'hFF;
ROM_MEM[10191] = 8'h2F;
ROM_MEM[10192] = 8'h11;
ROM_MEM[10193] = 8'h00;
ROM_MEM[10194] = 8'h00;
ROM_MEM[10195] = 8'h82;
ROM_MEM[10196] = 8'h09;
ROM_MEM[10197] = 8'h80;
ROM_MEM[10198] = 8'h48;
ROM_MEM[10199] = 8'h87;
ROM_MEM[10200] = 8'h03;
ROM_MEM[10201] = 8'h86;
ROM_MEM[10202] = 8'h01;
ROM_MEM[10203] = 8'h20;
ROM_MEM[10204] = 8'h40;
ROM_MEM[10205] = 8'h20;
ROM_MEM[10206] = 8'h40;
ROM_MEM[10207] = 8'h8E;
ROM_MEM[10208] = 8'h02;
ROM_MEM[10209] = 8'h20;
ROM_MEM[10210] = 8'h40;
ROM_MEM[10211] = 8'h1C;
ROM_MEM[10212] = 8'h30;
ROM_MEM[10213] = 8'h23;
ROM_MEM[10214] = 8'h10;
ROM_MEM[10215] = 8'h8F;
ROM_MEM[10216] = 8'h00;
ROM_MEM[10217] = 8'h20;
ROM_MEM[10218] = 8'h80;
ROM_MEM[10219] = 8'h20;
ROM_MEM[10220] = 8'h40;
ROM_MEM[10221] = 8'h20;
ROM_MEM[10222] = 8'h40;
ROM_MEM[10223] = 8'h20;
ROM_MEM[10224] = 8'h40;
ROM_MEM[10225] = 8'h1C;
ROM_MEM[10226] = 8'h30;
ROM_MEM[10227] = 8'h23;
ROM_MEM[10228] = 8'h10;
ROM_MEM[10229] = 8'h1F;
ROM_MEM[10230] = 8'h40;
ROM_MEM[10231] = 8'h1C;
ROM_MEM[10232] = 8'h30;
ROM_MEM[10233] = 8'h23;
ROM_MEM[10234] = 8'h10;
ROM_MEM[10235] = 8'h20;
ROM_MEM[10236] = 8'h60;
ROM_MEM[10237] = 8'h83;
ROM_MEM[10238] = 8'hFF;
ROM_MEM[10239] = 8'h20;
ROM_MEM[10240] = 8'h11;
ROM_MEM[10241] = 8'h83;
ROM_MEM[10242] = 8'hFF;
ROM_MEM[10243] = 8'h20;
ROM_MEM[10244] = 8'h11;
ROM_MEM[10245] = 8'h00;
ROM_MEM[10246] = 8'h00;
ROM_MEM[10247] = 8'h80;
ROM_MEM[10248] = 8'h3C;
ROM_MEM[10249] = 8'h90;
ROM_MEM[10250] = 8'h68;
ROM_MEM[10251] = 8'h39;
ROM_MEM[10252] = 8'h00;
ROM_MEM[10253] = 8'h00;
ROM_MEM[10254] = 8'h80;
ROM_MEM[10255] = 8'h3C;
ROM_MEM[10256] = 8'h8E;
ROM_MEM[10257] = 8'h02;
ROM_MEM[10258] = 8'h00;
ROM_MEM[10259] = 8'h40;
ROM_MEM[10260] = 8'h8F;
ROM_MEM[10261] = 8'h00;
ROM_MEM[10262] = 8'h85;
ROM_MEM[10263] = 8'h04;
ROM_MEM[10264] = 8'h90;
ROM_MEM[10265] = 8'h68;
ROM_MEM[10266] = 8'h39;
ROM_MEM[10267] = 8'h00;
ROM_MEM[10268] = 8'h00;
ROM_MEM[10269] = 8'h80;
ROM_MEM[10270] = 8'h3C;
ROM_MEM[10271] = 8'h8E;
ROM_MEM[10272] = 8'h04;
ROM_MEM[10273] = 8'h00;
ROM_MEM[10274] = 8'h40;
ROM_MEM[10275] = 8'h8F;
ROM_MEM[10276] = 8'h00;
ROM_MEM[10277] = 8'h90;
ROM_MEM[10278] = 8'h68;
ROM_MEM[10279] = 8'h48;
ROM_MEM[10280] = 8'h00;
ROM_MEM[10281] = 8'h00;
ROM_MEM[10282] = 8'h80;
ROM_MEM[10283] = 8'h3C;
ROM_MEM[10284] = 8'h8E;
ROM_MEM[10285] = 8'h06;
ROM_MEM[10286] = 8'h00;
ROM_MEM[10287] = 8'h40;
ROM_MEM[10288] = 8'h8F;
ROM_MEM[10289] = 8'h00;
ROM_MEM[10290] = 8'h85;
ROM_MEM[10291] = 8'h04;
ROM_MEM[10292] = 8'h90;
ROM_MEM[10293] = 8'h68;
ROM_MEM[10294] = 8'h48;
ROM_MEM[10295] = 8'h00;
ROM_MEM[10296] = 8'h00;
ROM_MEM[10297] = 8'h87;
ROM_MEM[10298] = 8'h01;
ROM_MEM[10299] = 8'h8E;
ROM_MEM[10300] = 8'h02;
ROM_MEM[10301] = 8'h31;
ROM_MEM[10302] = 8'h16;
ROM_MEM[10303] = 8'h31;
ROM_MEM[10304] = 8'h16;
ROM_MEM[10305] = 8'h31;
ROM_MEM[10306] = 8'h14;
ROM_MEM[10307] = 8'h85;
ROM_MEM[10308] = 8'h02;
ROM_MEM[10309] = 8'h8F;
ROM_MEM[10310] = 8'h00;
ROM_MEM[10311] = 8'h91;
ROM_MEM[10312] = 8'h87;
ROM_MEM[10313] = 8'h01;
ROM_MEM[10314] = 8'h8E;
ROM_MEM[10315] = 8'h02;
ROM_MEM[10316] = 8'h31;
ROM_MEM[10317] = 8'h10;
ROM_MEM[10318] = 8'h31;
ROM_MEM[10319] = 8'h10;
ROM_MEM[10320] = 8'h31;
ROM_MEM[10321] = 8'h10;
ROM_MEM[10322] = 8'h31;
ROM_MEM[10323] = 8'h10;
ROM_MEM[10324] = 8'h85;
ROM_MEM[10325] = 8'h02;
ROM_MEM[10326] = 8'h8F;
ROM_MEM[10327] = 8'h00;
ROM_MEM[10328] = 8'h91;
ROM_MEM[10329] = 8'h01;
ROM_MEM[10330] = 8'h02;
ROM_MEM[10331] = 8'h06;
ROM_MEM[10332] = 8'h00;
ROM_MEM[10333] = 8'h02;
ROM_MEM[10334] = 8'h02;
ROM_MEM[10335] = 8'h15;
ROM_MEM[10336] = 8'h04;
ROM_MEM[10337] = 8'h02;
ROM_MEM[10338] = 8'h02;
ROM_MEM[10339] = 8'h13;
ROM_MEM[10340] = 8'hF3;
ROM_MEM[10341] = 8'h01;
ROM_MEM[10342] = 8'h02;
ROM_MEM[10343] = 8'h11;
ROM_MEM[10344] = 8'h00;
ROM_MEM[10345] = 8'h01;
ROM_MEM[10346] = 8'h12;
ROM_MEM[10347] = 8'h01;
ROM_MEM[10348] = 8'h00;
ROM_MEM[10349] = 8'h15;
ROM_MEM[10350] = 8'h02;
ROM_MEM[10351] = 8'h09;
ROM_MEM[10352] = 8'h01;
ROM_MEM[10353] = 8'h01;
ROM_MEM[10354] = 8'h02;
ROM_MEM[10355] = 8'h1D;
ROM_MEM[10356] = 8'h00;
ROM_MEM[10357] = 8'h81;
ROM_MEM[10358] = 8'h02;
ROM_MEM[10359] = 8'h1F;
ROM_MEM[10360] = 8'h01;
ROM_MEM[10361] = 8'h04;
ROM_MEM[10362] = 8'h02;
ROM_MEM[10363] = 8'h21;
ROM_MEM[10364] = 8'h01;
ROM_MEM[10365] = 8'h02;
ROM_MEM[10366] = 8'h02;
ROM_MEM[10367] = 8'h26;
ROM_MEM[10368] = 8'h02;
ROM_MEM[10369] = 8'h01;
ROM_MEM[10370] = 8'h02;
ROM_MEM[10371] = 8'h2B;
ROM_MEM[10372] = 8'h00;
ROM_MEM[10373] = 8'h01;
ROM_MEM[10374] = 8'h10;
ROM_MEM[10375] = 8'h20;
ROM_MEM[10376] = 8'h00;
ROM_MEM[10377] = 8'h01;
ROM_MEM[10378] = 8'h06;
ROM_MEM[10379] = 8'h2B;
ROM_MEM[10380] = 8'h00;
ROM_MEM[10381] = 8'h02;
ROM_MEM[10382] = 8'h0A;
ROM_MEM[10383] = 8'h2A;
ROM_MEM[10384] = 8'hFF;
ROM_MEM[10385] = 8'h02;
ROM_MEM[10386] = 8'h0C;
ROM_MEM[10387] = 8'h28;
ROM_MEM[10388] = 8'hFF;
ROM_MEM[10389] = 8'h01;
ROM_MEM[10390] = 8'h0E;
ROM_MEM[10391] = 8'h26;
ROM_MEM[10392] = 8'h00;
ROM_MEM[10393] = 8'h01;
ROM_MEM[10394] = 8'h10;
ROM_MEM[10395] = 8'h25;
ROM_MEM[10396] = 8'h00;
ROM_MEM[10397] = 8'h01;
ROM_MEM[10398] = 8'h12;
ROM_MEM[10399] = 8'h24;
ROM_MEM[10400] = 8'h00;
ROM_MEM[10401] = 8'h01;
ROM_MEM[10402] = 8'h14;
ROM_MEM[10403] = 8'h23;
ROM_MEM[10404] = 8'h00;
ROM_MEM[10405] = 8'h01;
ROM_MEM[10406] = 8'h26;
ROM_MEM[10407] = 8'h22;
ROM_MEM[10408] = 8'h00;
ROM_MEM[10409] = 8'h01;
ROM_MEM[10410] = 8'h32;
ROM_MEM[10411] = 8'h21;
ROM_MEM[10412] = 8'h00;
ROM_MEM[10413] = 8'h00;
ROM_MEM[10414] = 8'h01;
ROM_MEM[10415] = 8'h12;
ROM_MEM[10416] = 8'h1B;
ROM_MEM[10417] = 8'h00;
ROM_MEM[10418] = 8'h02;
ROM_MEM[10419] = 8'h02;
ROM_MEM[10420] = 8'h15;
ROM_MEM[10421] = 8'h04;
ROM_MEM[10422] = 8'h02;
ROM_MEM[10423] = 8'h02;
ROM_MEM[10424] = 8'h0C;
ROM_MEM[10425] = 8'h05;
ROM_MEM[10426] = 8'h01;
ROM_MEM[10427] = 8'h02;
ROM_MEM[10428] = 8'h00;
ROM_MEM[10429] = 8'h00;
ROM_MEM[10430] = 8'h01;
ROM_MEM[10431] = 8'h12;
ROM_MEM[10432] = 8'h0A;
ROM_MEM[10433] = 8'h00;
ROM_MEM[10434] = 8'h14;
ROM_MEM[10435] = 8'h02;
ROM_MEM[10436] = 8'h0A;
ROM_MEM[10437] = 8'h01;
ROM_MEM[10438] = 8'h01;
ROM_MEM[10439] = 8'h02;
ROM_MEM[10440] = 8'h1D;
ROM_MEM[10441] = 8'h00;
ROM_MEM[10442] = 8'h2B;
ROM_MEM[10443] = 8'h02;
ROM_MEM[10444] = 8'h1F;
ROM_MEM[10445] = 8'h01;
ROM_MEM[10446] = 8'h08;
ROM_MEM[10447] = 8'h02;
ROM_MEM[10448] = 8'h37;
ROM_MEM[10449] = 8'hFF;
ROM_MEM[10450] = 8'h6D;
ROM_MEM[10451] = 8'h02;
ROM_MEM[10452] = 8'h1F;
ROM_MEM[10453] = 8'h01;
ROM_MEM[10454] = 8'h01;
ROM_MEM[10455] = 8'h10;
ROM_MEM[10456] = 8'h40;
ROM_MEM[10457] = 8'h00;
ROM_MEM[10458] = 8'h06;
ROM_MEM[10459] = 8'h02;
ROM_MEM[10460] = 8'h41;
ROM_MEM[10461] = 8'h02;
ROM_MEM[10462] = 8'h01;
ROM_MEM[10463] = 8'h12;
ROM_MEM[10464] = 8'h40;
ROM_MEM[10465] = 8'h00;
ROM_MEM[10466] = 8'h03;
ROM_MEM[10467] = 8'h08;
ROM_MEM[10468] = 8'h8B;
ROM_MEM[10469] = 8'hFF;
ROM_MEM[10470] = 8'h02;
ROM_MEM[10471] = 8'h0A;
ROM_MEM[10472] = 8'h88;
ROM_MEM[10473] = 8'hFF;
ROM_MEM[10474] = 8'h01;
ROM_MEM[10475] = 8'h0C;
ROM_MEM[10476] = 8'h86;
ROM_MEM[10477] = 8'h00;
ROM_MEM[10478] = 8'h01;
ROM_MEM[10479] = 8'h0E;
ROM_MEM[10480] = 8'h85;
ROM_MEM[10481] = 8'h00;
ROM_MEM[10482] = 8'h01;
ROM_MEM[10483] = 8'h16;
ROM_MEM[10484] = 8'h84;
ROM_MEM[10485] = 8'h00;
ROM_MEM[10486] = 8'h01;
ROM_MEM[10487] = 8'hD0;
ROM_MEM[10488] = 8'h83;
ROM_MEM[10489] = 8'h00;
ROM_MEM[10490] = 8'h01;
ROM_MEM[10491] = 8'h22;
ROM_MEM[10492] = 8'h82;
ROM_MEM[10493] = 8'h00;
ROM_MEM[10494] = 8'h01;
ROM_MEM[10495] = 8'h1C;
ROM_MEM[10496] = 8'h81;
ROM_MEM[10497] = 8'h00;
ROM_MEM[10498] = 8'h00;
ROM_MEM[10499] = 8'h03;
ROM_MEM[10500] = 8'h0A;
ROM_MEM[10501] = 8'h0C;
ROM_MEM[10502] = 8'h01;
ROM_MEM[10503] = 8'h02;
ROM_MEM[10504] = 8'h08;
ROM_MEM[10505] = 8'h0F;
ROM_MEM[10506] = 8'h01;
ROM_MEM[10507] = 8'h01;
ROM_MEM[10508] = 8'h06;
ROM_MEM[10509] = 8'h11;
ROM_MEM[10510] = 8'h00;
ROM_MEM[10511] = 8'h01;
ROM_MEM[10512] = 8'h06;
ROM_MEM[10513] = 8'h12;
ROM_MEM[10514] = 8'h00;
ROM_MEM[10515] = 8'h03;
ROM_MEM[10516] = 8'h04;
ROM_MEM[10517] = 8'h11;
ROM_MEM[10518] = 8'hFF;
ROM_MEM[10519] = 8'h06;
ROM_MEM[10520] = 8'h02;
ROM_MEM[10521] = 8'h0E;
ROM_MEM[10522] = 8'hFF;
ROM_MEM[10523] = 8'h3B;
ROM_MEM[10524] = 8'h02;
ROM_MEM[10525] = 8'h0A;
ROM_MEM[10526] = 8'h01;
ROM_MEM[10527] = 8'h01;
ROM_MEM[10528] = 8'h1A;
ROM_MEM[10529] = 8'h81;
ROM_MEM[10530] = 8'h00;
ROM_MEM[10531] = 8'h01;
ROM_MEM[10532] = 8'h10;
ROM_MEM[10533] = 8'h82;
ROM_MEM[10534] = 8'h00;
ROM_MEM[10535] = 8'h01;
ROM_MEM[10536] = 8'h06;
ROM_MEM[10537] = 8'h83;
ROM_MEM[10538] = 8'h00;
ROM_MEM[10539] = 8'h01;
ROM_MEM[10540] = 8'h04;
ROM_MEM[10541] = 8'h84;
ROM_MEM[10542] = 8'h00;
ROM_MEM[10543] = 8'h01;
ROM_MEM[10544] = 8'h06;
ROM_MEM[10545] = 8'h85;
ROM_MEM[10546] = 8'h00;
ROM_MEM[10547] = 8'h02;
ROM_MEM[10548] = 8'h04;
ROM_MEM[10549] = 8'h86;
ROM_MEM[10550] = 8'h01;
ROM_MEM[10551] = 8'h08;
ROM_MEM[10552] = 8'h02;
ROM_MEM[10553] = 8'h88;
ROM_MEM[10554] = 8'h01;
ROM_MEM[10555] = 8'h01;
ROM_MEM[10556] = 8'h02;
ROM_MEM[10557] = 8'h8F;
ROM_MEM[10558] = 8'h00;
ROM_MEM[10559] = 8'h01;
ROM_MEM[10560] = 8'h04;
ROM_MEM[10561] = 8'h8E;
ROM_MEM[10562] = 8'h00;
ROM_MEM[10563] = 8'h01;
ROM_MEM[10564] = 8'h06;
ROM_MEM[10565] = 8'h8D;
ROM_MEM[10566] = 8'h00;
ROM_MEM[10567] = 8'h02;
ROM_MEM[10568] = 8'h04;
ROM_MEM[10569] = 8'h8C;
ROM_MEM[10570] = 8'hFF;
ROM_MEM[10571] = 8'h02;
ROM_MEM[10572] = 8'h06;
ROM_MEM[10573] = 8'h8A;
ROM_MEM[10574] = 8'hFF;
ROM_MEM[10575] = 8'h07;
ROM_MEM[10576] = 8'h08;
ROM_MEM[10577] = 8'h88;
ROM_MEM[10578] = 8'hFF;
ROM_MEM[10579] = 8'h01;
ROM_MEM[10580] = 8'h1C;
ROM_MEM[10581] = 8'h81;
ROM_MEM[10582] = 8'h00;
ROM_MEM[10583] = 8'h00;
ROM_MEM[10584] = 8'h02;
ROM_MEM[10585] = 8'h02;
ROM_MEM[10586] = 8'h81;
ROM_MEM[10587] = 8'h01;
ROM_MEM[10588] = 8'h02;
ROM_MEM[10589] = 8'h02;
ROM_MEM[10590] = 8'h84;
ROM_MEM[10591] = 8'h03;
ROM_MEM[10592] = 8'h01;
ROM_MEM[10593] = 8'h02;
ROM_MEM[10594] = 8'h8B;
ROM_MEM[10595] = 8'h00;
ROM_MEM[10596] = 8'h02;
ROM_MEM[10597] = 8'h04;
ROM_MEM[10598] = 8'h8F;
ROM_MEM[10599] = 8'hFF;
ROM_MEM[10600] = 8'h01;
ROM_MEM[10601] = 8'h06;
ROM_MEM[10602] = 8'h8D;
ROM_MEM[10603] = 8'h00;
ROM_MEM[10604] = 8'h02;
ROM_MEM[10605] = 8'h04;
ROM_MEM[10606] = 8'h8C;
ROM_MEM[10607] = 8'hFF;
ROM_MEM[10608] = 8'h02;
ROM_MEM[10609] = 8'h06;
ROM_MEM[10610] = 8'h8A;
ROM_MEM[10611] = 8'hFF;
ROM_MEM[10612] = 8'h07;
ROM_MEM[10613] = 8'h08;
ROM_MEM[10614] = 8'h88;
ROM_MEM[10615] = 8'hFF;
ROM_MEM[10616] = 8'h01;
ROM_MEM[10617] = 8'h1C;
ROM_MEM[10618] = 8'h81;
ROM_MEM[10619] = 8'h00;
ROM_MEM[10620] = 8'h00;
ROM_MEM[10621] = 8'h01;
ROM_MEM[10622] = 8'h34;
ROM_MEM[10623] = 8'h23;
ROM_MEM[10624] = 8'h00;
ROM_MEM[10625] = 8'h09;
ROM_MEM[10626] = 8'h02;
ROM_MEM[10627] = 8'h23;
ROM_MEM[10628] = 8'hFF;
ROM_MEM[10629] = 8'h06;
ROM_MEM[10630] = 8'h02;
ROM_MEM[10631] = 8'h1A;
ROM_MEM[10632] = 8'hFF;
ROM_MEM[10633] = 8'h17;
ROM_MEM[10634] = 8'h02;
ROM_MEM[10635] = 8'h16;
ROM_MEM[10636] = 8'h01;
ROM_MEM[10637] = 8'h01;
ROM_MEM[10638] = 8'h34;
ROM_MEM[10639] = 8'hC0;
ROM_MEM[10640] = 8'h00;
ROM_MEM[10641] = 8'h0F;
ROM_MEM[10642] = 8'h02;
ROM_MEM[10643] = 8'hC1;
ROM_MEM[10644] = 8'h01;
ROM_MEM[10645] = 8'h01;
ROM_MEM[10646] = 8'h02;
ROM_MEM[10647] = 8'hCF;
ROM_MEM[10648] = 8'h00;
ROM_MEM[10649] = 8'h02;
ROM_MEM[10650] = 8'h04;
ROM_MEM[10651] = 8'hCE;
ROM_MEM[10652] = 8'hFF;
ROM_MEM[10653] = 8'h01;
ROM_MEM[10654] = 8'h02;
ROM_MEM[10655] = 8'hCC;
ROM_MEM[10656] = 8'h00;
ROM_MEM[10657] = 8'h01;
ROM_MEM[10658] = 8'h04;
ROM_MEM[10659] = 8'hCB;
ROM_MEM[10660] = 8'h00;
ROM_MEM[10661] = 8'h01;
ROM_MEM[10662] = 8'h02;
ROM_MEM[10663] = 8'hCA;
ROM_MEM[10664] = 8'h00;
ROM_MEM[10665] = 8'h01;
ROM_MEM[10666] = 8'h04;
ROM_MEM[10667] = 8'hC9;
ROM_MEM[10668] = 8'h00;
ROM_MEM[10669] = 8'h01;
ROM_MEM[10670] = 8'h02;
ROM_MEM[10671] = 8'hC8;
ROM_MEM[10672] = 8'h00;
ROM_MEM[10673] = 8'h01;
ROM_MEM[10674] = 8'h04;
ROM_MEM[10675] = 8'hC7;
ROM_MEM[10676] = 8'h00;
ROM_MEM[10677] = 8'h05;
ROM_MEM[10678] = 8'h02;
ROM_MEM[10679] = 8'hC6;
ROM_MEM[10680] = 8'hFF;
ROM_MEM[10681] = 8'h01;
ROM_MEM[10682] = 8'h02;
ROM_MEM[10683] = 8'hC2;
ROM_MEM[10684] = 8'h00;
ROM_MEM[10685] = 8'h01;
ROM_MEM[10686] = 8'h04;
ROM_MEM[10687] = 8'hC1;
ROM_MEM[10688] = 8'h00;
ROM_MEM[10689] = 8'h00;
ROM_MEM[10690] = 8'h02;
ROM_MEM[10691] = 8'h02;
ROM_MEM[10692] = 8'hC1;
ROM_MEM[10693] = 8'h01;
ROM_MEM[10694] = 8'h02;
ROM_MEM[10695] = 8'h02;
ROM_MEM[10696] = 8'hC4;
ROM_MEM[10697] = 8'h03;
ROM_MEM[10698] = 8'h01;
ROM_MEM[10699] = 8'h02;
ROM_MEM[10700] = 8'hCB;
ROM_MEM[10701] = 8'h00;
ROM_MEM[10702] = 8'h03;
ROM_MEM[10703] = 8'h04;
ROM_MEM[10704] = 8'hCF;
ROM_MEM[10705] = 8'hFF;
ROM_MEM[10706] = 8'h01;
ROM_MEM[10707] = 8'h02;
ROM_MEM[10708] = 8'hCC;
ROM_MEM[10709] = 8'h00;
ROM_MEM[10710] = 8'h01;
ROM_MEM[10711] = 8'h04;
ROM_MEM[10712] = 8'hCB;
ROM_MEM[10713] = 8'h00;
ROM_MEM[10714] = 8'h01;
ROM_MEM[10715] = 8'h02;
ROM_MEM[10716] = 8'hCA;
ROM_MEM[10717] = 8'h00;
ROM_MEM[10718] = 8'h01;
ROM_MEM[10719] = 8'h04;
ROM_MEM[10720] = 8'hC9;
ROM_MEM[10721] = 8'h00;
ROM_MEM[10722] = 8'h01;
ROM_MEM[10723] = 8'h02;
ROM_MEM[10724] = 8'hC8;
ROM_MEM[10725] = 8'h00;
ROM_MEM[10726] = 8'h01;
ROM_MEM[10727] = 8'h04;
ROM_MEM[10728] = 8'hC7;
ROM_MEM[10729] = 8'h00;
ROM_MEM[10730] = 8'h04;
ROM_MEM[10731] = 8'h02;
ROM_MEM[10732] = 8'hC6;
ROM_MEM[10733] = 8'h00;
ROM_MEM[10734] = 8'h02;
ROM_MEM[10735] = 8'h04;
ROM_MEM[10736] = 8'hC2;
ROM_MEM[10737] = 8'hFF;
ROM_MEM[10738] = 8'h00;
ROM_MEM[10739] = 8'h01;
ROM_MEM[10740] = 8'h38;
ROM_MEM[10741] = 8'h03;
ROM_MEM[10742] = 8'h00;
ROM_MEM[10743] = 8'h01;
ROM_MEM[10744] = 8'h0A;
ROM_MEM[10745] = 8'h41;
ROM_MEM[10746] = 8'h00;
ROM_MEM[10747] = 8'h01;
ROM_MEM[10748] = 8'h08;
ROM_MEM[10749] = 8'h42;
ROM_MEM[10750] = 8'h00;
ROM_MEM[10751] = 8'h01;
ROM_MEM[10752] = 8'h06;
ROM_MEM[10753] = 8'h43;
ROM_MEM[10754] = 8'h00;
ROM_MEM[10755] = 8'h01;
ROM_MEM[10756] = 8'h04;
ROM_MEM[10757] = 8'h44;
ROM_MEM[10758] = 8'h00;
ROM_MEM[10759] = 8'h08;
ROM_MEM[10760] = 8'h02;
ROM_MEM[10761] = 8'h45;
ROM_MEM[10762] = 8'h01;
ROM_MEM[10763] = 8'h02;
ROM_MEM[10764] = 8'h01;
ROM_MEM[10765] = 8'h4D;
ROM_MEM[10766] = 8'h01;
ROM_MEM[10767] = 8'h01;
ROM_MEM[10768] = 8'h0A;
ROM_MEM[10769] = 8'h4F;
ROM_MEM[10770] = 8'h00;
ROM_MEM[10771] = 8'h00;
ROM_MEM[10772] = 8'h08;
ROM_MEM[10773] = 8'h02;
ROM_MEM[10774] = 8'h56;
ROM_MEM[10775] = 8'hF8;
ROM_MEM[10776] = 8'h03;
ROM_MEM[10777] = 8'h02;
ROM_MEM[10778] = 8'h81;
ROM_MEM[10779] = 8'h01;
ROM_MEM[10780] = 8'h02;
ROM_MEM[10781] = 8'h02;
ROM_MEM[10782] = 8'h86;
ROM_MEM[10783] = 8'h04;
ROM_MEM[10784] = 8'h03;
ROM_MEM[10785] = 8'h02;
ROM_MEM[10786] = 8'h8C;
ROM_MEM[10787] = 8'h01;
ROM_MEM[10788] = 8'h00;
ROM_MEM[10789] = 8'h02;
ROM_MEM[10790] = 8'h02;
ROM_MEM[10791] = 8'h23;
ROM_MEM[10792] = 8'hFF;
ROM_MEM[10793] = 8'h01;
ROM_MEM[10794] = 8'h0A;
ROM_MEM[10795] = 8'h22;
ROM_MEM[10796] = 8'h00;
ROM_MEM[10797] = 8'h2F;
ROM_MEM[10798] = 8'h02;
ROM_MEM[10799] = 8'h02;
ROM_MEM[10800] = 8'h01;
ROM_MEM[10801] = 8'h01;
ROM_MEM[10802] = 8'h04;
ROM_MEM[10803] = 8'h2F;
ROM_MEM[10804] = 8'h00;
ROM_MEM[10805] = 8'h01;
ROM_MEM[10806] = 8'h0A;
ROM_MEM[10807] = 8'h20;
ROM_MEM[10808] = 8'h00;
ROM_MEM[10809] = 8'h03;
ROM_MEM[10810] = 8'h02;
ROM_MEM[10811] = 8'h2F;
ROM_MEM[10812] = 8'hFF;
ROM_MEM[10813] = 8'h03;
ROM_MEM[10814] = 8'h04;
ROM_MEM[10815] = 8'h2C;
ROM_MEM[10816] = 8'hFF;
ROM_MEM[10817] = 8'h03;
ROM_MEM[10818] = 8'h06;
ROM_MEM[10819] = 8'h29;
ROM_MEM[10820] = 8'hFF;
ROM_MEM[10821] = 8'h02;
ROM_MEM[10822] = 8'h08;
ROM_MEM[10823] = 8'h26;
ROM_MEM[10824] = 8'hFF;
ROM_MEM[10825] = 8'h01;
ROM_MEM[10826] = 8'h04;
ROM_MEM[10827] = 8'h24;
ROM_MEM[10828] = 8'h00;
ROM_MEM[10829] = 8'h02;
ROM_MEM[10830] = 8'h02;
ROM_MEM[10831] = 8'h04;
ROM_MEM[10832] = 8'h20;
ROM_MEM[10833] = 8'h02;
ROM_MEM[10834] = 8'h0A;
ROM_MEM[10835] = 8'h23;
ROM_MEM[10836] = 8'hFF;
ROM_MEM[10837] = 8'h01;
ROM_MEM[10838] = 8'h0C;
ROM_MEM[10839] = 8'h21;
ROM_MEM[10840] = 8'h00;
ROM_MEM[10841] = 8'h00;
ROM_MEM[10842] = 8'h05;
ROM_MEM[10843] = 8'h02;
ROM_MEM[10844] = 8'h16;
ROM_MEM[10845] = 8'h01;
ROM_MEM[10846] = 8'h03;
ROM_MEM[10847] = 8'h02;
ROM_MEM[10848] = 8'h19;
ROM_MEM[10849] = 8'hFF;
ROM_MEM[10850] = 8'h05;
ROM_MEM[10851] = 8'h02;
ROM_MEM[10852] = 8'h16;
ROM_MEM[10853] = 8'h01;
ROM_MEM[10854] = 8'h03;
ROM_MEM[10855] = 8'h02;
ROM_MEM[10856] = 8'h19;
ROM_MEM[10857] = 8'hFF;
ROM_MEM[10858] = 8'h05;
ROM_MEM[10859] = 8'h02;
ROM_MEM[10860] = 8'h16;
ROM_MEM[10861] = 8'h01;
ROM_MEM[10862] = 8'h03;
ROM_MEM[10863] = 8'h02;
ROM_MEM[10864] = 8'h19;
ROM_MEM[10865] = 8'hFF;
ROM_MEM[10866] = 8'h05;
ROM_MEM[10867] = 8'h02;
ROM_MEM[10868] = 8'h16;
ROM_MEM[10869] = 8'h01;
ROM_MEM[10870] = 8'h03;
ROM_MEM[10871] = 8'h02;
ROM_MEM[10872] = 8'h19;
ROM_MEM[10873] = 8'hFF;
ROM_MEM[10874] = 8'h05;
ROM_MEM[10875] = 8'h02;
ROM_MEM[10876] = 8'h16;
ROM_MEM[10877] = 8'h01;
ROM_MEM[10878] = 8'h03;
ROM_MEM[10879] = 8'h02;
ROM_MEM[10880] = 8'h19;
ROM_MEM[10881] = 8'hFF;
ROM_MEM[10882] = 8'h05;
ROM_MEM[10883] = 8'h02;
ROM_MEM[10884] = 8'h16;
ROM_MEM[10885] = 8'h01;
ROM_MEM[10886] = 8'h03;
ROM_MEM[10887] = 8'h02;
ROM_MEM[10888] = 8'h19;
ROM_MEM[10889] = 8'hFF;
ROM_MEM[10890] = 8'h03;
ROM_MEM[10891] = 8'h02;
ROM_MEM[10892] = 8'h16;
ROM_MEM[10893] = 8'h01;
ROM_MEM[10894] = 8'h01;
ROM_MEM[10895] = 8'h04;
ROM_MEM[10896] = 8'h0F;
ROM_MEM[10897] = 8'h00;
ROM_MEM[10898] = 8'h01;
ROM_MEM[10899] = 8'h06;
ROM_MEM[10900] = 8'h00;
ROM_MEM[10901] = 8'h00;
ROM_MEM[10902] = 8'h03;
ROM_MEM[10903] = 8'h0A;
ROM_MEM[10904] = 8'h0F;
ROM_MEM[10905] = 8'hFF;
ROM_MEM[10906] = 8'h09;
ROM_MEM[10907] = 8'h04;
ROM_MEM[10908] = 8'h0C;
ROM_MEM[10909] = 8'hFF;
ROM_MEM[10910] = 8'h01;
ROM_MEM[10911] = 8'h06;
ROM_MEM[10912] = 8'h03;
ROM_MEM[10913] = 8'h00;
ROM_MEM[10914] = 8'h01;
ROM_MEM[10915] = 8'h08;
ROM_MEM[10916] = 8'h02;
ROM_MEM[10917] = 8'h00;
ROM_MEM[10918] = 8'h01;
ROM_MEM[10919] = 8'h0C;
ROM_MEM[10920] = 8'h01;
ROM_MEM[10921] = 8'h00;
ROM_MEM[10922] = 8'h00;
ROM_MEM[10923] = 8'h02;
ROM_MEM[10924] = 8'h90;
ROM_MEM[10925] = 8'h46;
ROM_MEM[10926] = 8'h00;
ROM_MEM[10927] = 8'h02;
ROM_MEM[10928] = 8'h90;
ROM_MEM[10929] = 8'h47;
ROM_MEM[10930] = 8'h00;
ROM_MEM[10931] = 8'h02;
ROM_MEM[10932] = 8'h90;
ROM_MEM[10933] = 8'h48;
ROM_MEM[10934] = 8'h00;
ROM_MEM[10935] = 8'h02;
ROM_MEM[10936] = 8'h90;
ROM_MEM[10937] = 8'h49;
ROM_MEM[10938] = 8'h00;
ROM_MEM[10939] = 8'h02;
ROM_MEM[10940] = 8'h90;
ROM_MEM[10941] = 8'h4B;
ROM_MEM[10942] = 8'h00;
ROM_MEM[10943] = 8'h02;
ROM_MEM[10944] = 8'h90;
ROM_MEM[10945] = 8'h4C;
ROM_MEM[10946] = 8'h00;
ROM_MEM[10947] = 8'h02;
ROM_MEM[10948] = 8'h90;
ROM_MEM[10949] = 8'h4D;
ROM_MEM[10950] = 8'h00;
ROM_MEM[10951] = 8'h02;
ROM_MEM[10952] = 8'h90;
ROM_MEM[10953] = 8'h4E;
ROM_MEM[10954] = 8'h00;
ROM_MEM[10955] = 8'h01;
ROM_MEM[10956] = 8'h0A;
ROM_MEM[10957] = 8'h4F;
ROM_MEM[10958] = 8'h00;
ROM_MEM[10959] = 8'h01;
ROM_MEM[10960] = 8'h08;
ROM_MEM[10961] = 8'h40;
ROM_MEM[10962] = 8'h00;
ROM_MEM[10963] = 8'h01;
ROM_MEM[10964] = 8'h04;
ROM_MEM[10965] = 8'h4F;
ROM_MEM[10966] = 8'h00;
ROM_MEM[10967] = 8'h01;
ROM_MEM[10968] = 8'h06;
ROM_MEM[10969] = 8'h4E;
ROM_MEM[10970] = 8'h00;
ROM_MEM[10971] = 8'h01;
ROM_MEM[10972] = 8'h08;
ROM_MEM[10973] = 8'h4D;
ROM_MEM[10974] = 8'h00;
ROM_MEM[10975] = 8'h01;
ROM_MEM[10976] = 8'h0A;
ROM_MEM[10977] = 8'h4C;
ROM_MEM[10978] = 8'h00;
ROM_MEM[10979] = 8'h01;
ROM_MEM[10980] = 8'h0C;
ROM_MEM[10981] = 8'h4B;
ROM_MEM[10982] = 8'h00;
ROM_MEM[10983] = 8'h01;
ROM_MEM[10984] = 8'h0E;
ROM_MEM[10985] = 8'h4A;
ROM_MEM[10986] = 8'h00;
ROM_MEM[10987] = 8'h01;
ROM_MEM[10988] = 8'h10;
ROM_MEM[10989] = 8'h49;
ROM_MEM[10990] = 8'h00;
ROM_MEM[10991] = 8'h01;
ROM_MEM[10992] = 8'h12;
ROM_MEM[10993] = 8'h48;
ROM_MEM[10994] = 8'h00;
ROM_MEM[10995] = 8'h01;
ROM_MEM[10996] = 8'h14;
ROM_MEM[10997] = 8'h47;
ROM_MEM[10998] = 8'h00;
ROM_MEM[10999] = 8'h01;
ROM_MEM[11000] = 8'h16;
ROM_MEM[11001] = 8'h46;
ROM_MEM[11002] = 8'h00;
ROM_MEM[11003] = 8'h01;
ROM_MEM[11004] = 8'h18;
ROM_MEM[11005] = 8'h45;
ROM_MEM[11006] = 8'h00;
ROM_MEM[11007] = 8'h01;
ROM_MEM[11008] = 8'h1A;
ROM_MEM[11009] = 8'h44;
ROM_MEM[11010] = 8'h00;
ROM_MEM[11011] = 8'h01;
ROM_MEM[11012] = 8'h1C;
ROM_MEM[11013] = 8'h43;
ROM_MEM[11014] = 8'h00;
ROM_MEM[11015] = 8'h01;
ROM_MEM[11016] = 8'h1E;
ROM_MEM[11017] = 8'h42;
ROM_MEM[11018] = 8'h00;
ROM_MEM[11019] = 8'h01;
ROM_MEM[11020] = 8'h20;
ROM_MEM[11021] = 8'h41;
ROM_MEM[11022] = 8'h00;
ROM_MEM[11023] = 8'h00;
ROM_MEM[11024] = 8'h01;
ROM_MEM[11025] = 8'h5A;
ROM_MEM[11026] = 8'h41;
ROM_MEM[11027] = 8'h00;
ROM_MEM[11028] = 8'h01;
ROM_MEM[11029] = 8'h5A;
ROM_MEM[11030] = 8'h3E;
ROM_MEM[11031] = 8'h00;
ROM_MEM[11032] = 8'h01;
ROM_MEM[11033] = 8'h1A;
ROM_MEM[11034] = 8'h4F;
ROM_MEM[11035] = 8'h00;
ROM_MEM[11036] = 8'h02;
ROM_MEM[11037] = 8'h02;
ROM_MEM[11038] = 8'h4E;
ROM_MEM[11039] = 8'hFF;
ROM_MEM[11040] = 8'h09;
ROM_MEM[11041] = 8'h04;
ROM_MEM[11042] = 8'h4C;
ROM_MEM[11043] = 8'hFF;
ROM_MEM[11044] = 8'h01;
ROM_MEM[11045] = 8'h06;
ROM_MEM[11046] = 8'h43;
ROM_MEM[11047] = 8'h00;
ROM_MEM[11048] = 8'h01;
ROM_MEM[11049] = 8'h08;
ROM_MEM[11050] = 8'h42;
ROM_MEM[11051] = 8'h00;
ROM_MEM[11052] = 8'h01;
ROM_MEM[11053] = 8'h0A;
ROM_MEM[11054] = 8'h41;
ROM_MEM[11055] = 8'h00;
ROM_MEM[11056] = 8'h00;
ROM_MEM[11057] = 8'h01;
ROM_MEM[11058] = 8'h0E;
ROM_MEM[11059] = 8'h08;
ROM_MEM[11060] = 8'h00;
ROM_MEM[11061] = 8'h01;
ROM_MEM[11062] = 8'h02;
ROM_MEM[11063] = 8'h41;
ROM_MEM[11064] = 8'h00;
ROM_MEM[11065] = 8'h07;
ROM_MEM[11066] = 8'h01;
ROM_MEM[11067] = 8'h42;
ROM_MEM[11068] = 8'h01;
ROM_MEM[11069] = 8'h03;
ROM_MEM[11070] = 8'h01;
ROM_MEM[11071] = 8'h4A;
ROM_MEM[11072] = 8'h02;
ROM_MEM[11073] = 8'h01;
ROM_MEM[11074] = 8'h02;
ROM_MEM[11075] = 8'h4F;
ROM_MEM[11076] = 8'h00;
ROM_MEM[11077] = 8'h00;
ROM_MEM[11078] = 8'h32;
ROM_MEM[11079] = 8'h01;
ROM_MEM[11080] = 8'h37;
ROM_MEM[11081] = 8'h04;
ROM_MEM[11082] = 8'h01;
ROM_MEM[11083] = 8'h02;
ROM_MEM[11084] = 8'hFF;
ROM_MEM[11085] = 8'h00;
ROM_MEM[11086] = 8'h01;
ROM_MEM[11087] = 8'h0C;
ROM_MEM[11088] = 8'hA9;
ROM_MEM[11089] = 8'h00;
ROM_MEM[11090] = 8'h01;
ROM_MEM[11091] = 8'h0A;
ROM_MEM[11092] = 8'hA8;
ROM_MEM[11093] = 8'h00;
ROM_MEM[11094] = 8'h01;
ROM_MEM[11095] = 8'h08;
ROM_MEM[11096] = 8'hA7;
ROM_MEM[11097] = 8'h00;
ROM_MEM[11098] = 8'h01;
ROM_MEM[11099] = 8'h06;
ROM_MEM[11100] = 8'hA6;
ROM_MEM[11101] = 8'h00;
ROM_MEM[11102] = 8'h01;
ROM_MEM[11103] = 8'h04;
ROM_MEM[11104] = 8'hA5;
ROM_MEM[11105] = 8'h00;
ROM_MEM[11106] = 8'h05;
ROM_MEM[11107] = 8'h02;
ROM_MEM[11108] = 8'hA4;
ROM_MEM[11109] = 8'hFF;
ROM_MEM[11110] = 8'h01;
ROM_MEM[11111] = 8'h02;
ROM_MEM[11112] = 8'hA1;
ROM_MEM[11113] = 8'h00;
ROM_MEM[11114] = 8'h00;
ROM_MEM[11115] = 8'h01;
ROM_MEM[11116] = 8'h08;
ROM_MEM[11117] = 8'h05;
ROM_MEM[11118] = 8'h00;
ROM_MEM[11119] = 8'h2C;
ROM_MEM[11120] = 8'h01;
ROM_MEM[11121] = 8'h37;
ROM_MEM[11122] = 8'h04;
ROM_MEM[11123] = 8'h01;
ROM_MEM[11124] = 8'h08;
ROM_MEM[11125] = 8'h47;
ROM_MEM[11126] = 8'h00;
ROM_MEM[11127] = 8'h01;
ROM_MEM[11128] = 8'h16;
ROM_MEM[11129] = 8'hA7;
ROM_MEM[11130] = 8'h00;
ROM_MEM[11131] = 8'h01;
ROM_MEM[11132] = 8'h06;
ROM_MEM[11133] = 8'hA6;
ROM_MEM[11134] = 8'h00;
ROM_MEM[11135] = 8'h01;
ROM_MEM[11136] = 8'h04;
ROM_MEM[11137] = 8'hA5;
ROM_MEM[11138] = 8'h00;
ROM_MEM[11139] = 8'h05;
ROM_MEM[11140] = 8'h02;
ROM_MEM[11141] = 8'hA4;
ROM_MEM[11142] = 8'hFF;
ROM_MEM[11143] = 8'h01;
ROM_MEM[11144] = 8'h02;
ROM_MEM[11145] = 8'hA1;
ROM_MEM[11146] = 8'h00;
ROM_MEM[11147] = 8'h00;
ROM_MEM[11148] = 8'h05;
ROM_MEM[11149] = 8'h01;
ROM_MEM[11150] = 8'h23;
ROM_MEM[11151] = 8'h01;
ROM_MEM[11152] = 8'h0D;
ROM_MEM[11153] = 8'h01;
ROM_MEM[11154] = 8'h2A;
ROM_MEM[11155] = 8'h02;
ROM_MEM[11156] = 8'h09;
ROM_MEM[11157] = 8'h01;
ROM_MEM[11158] = 8'h45;
ROM_MEM[11159] = 8'h03;
ROM_MEM[11160] = 8'h08;
ROM_MEM[11161] = 8'h01;
ROM_MEM[11162] = 8'h61;
ROM_MEM[11163] = 8'h04;
ROM_MEM[11164] = 8'h04;
ROM_MEM[11165] = 8'h01;
ROM_MEM[11166] = 8'h83;
ROM_MEM[11167] = 8'h05;
ROM_MEM[11168] = 8'h05;
ROM_MEM[11169] = 8'h01;
ROM_MEM[11170] = 8'h99;
ROM_MEM[11171] = 8'h06;
ROM_MEM[11172] = 8'h04;
ROM_MEM[11173] = 8'h01;
ROM_MEM[11174] = 8'hB8;
ROM_MEM[11175] = 8'h07;
ROM_MEM[11176] = 8'h04;
ROM_MEM[11177] = 8'h01;
ROM_MEM[11178] = 8'hD5;
ROM_MEM[11179] = 8'h09;
ROM_MEM[11180] = 8'h11;
ROM_MEM[11181] = 8'h01;
ROM_MEM[11182] = 8'h2D;
ROM_MEM[11183] = 8'h02;
ROM_MEM[11184] = 8'h0A;
ROM_MEM[11185] = 8'h01;
ROM_MEM[11186] = 8'h4F;
ROM_MEM[11187] = 8'h03;
ROM_MEM[11188] = 8'h08;
ROM_MEM[11189] = 8'h01;
ROM_MEM[11190] = 8'h6E;
ROM_MEM[11191] = 8'h04;
ROM_MEM[11192] = 8'h05;
ROM_MEM[11193] = 8'h01;
ROM_MEM[11194] = 8'h90;
ROM_MEM[11195] = 8'h05;
ROM_MEM[11196] = 8'h07;
ROM_MEM[11197] = 8'h01;
ROM_MEM[11198] = 8'hAA;
ROM_MEM[11199] = 8'h06;
ROM_MEM[11200] = 8'h03;
ROM_MEM[11201] = 8'h01;
ROM_MEM[11202] = 8'hD7;
ROM_MEM[11203] = 8'h07;
ROM_MEM[11204] = 8'h02;
ROM_MEM[11205] = 8'h01;
ROM_MEM[11206] = 8'hED;
ROM_MEM[11207] = 8'h08;
ROM_MEM[11208] = 8'h04;
ROM_MEM[11209] = 8'h01;
ROM_MEM[11210] = 8'h33;
ROM_MEM[11211] = 8'h01;
ROM_MEM[11212] = 8'h09;
ROM_MEM[11213] = 8'h01;
ROM_MEM[11214] = 8'h38;
ROM_MEM[11215] = 8'h02;
ROM_MEM[11216] = 8'h0C;
ROM_MEM[11217] = 8'h01;
ROM_MEM[11218] = 8'h4B;
ROM_MEM[11219] = 8'h03;
ROM_MEM[11220] = 8'h07;
ROM_MEM[11221] = 8'h01;
ROM_MEM[11222] = 8'h6E;
ROM_MEM[11223] = 8'h04;
ROM_MEM[11224] = 8'h08;
ROM_MEM[11225] = 8'h01;
ROM_MEM[11226] = 8'h8A;
ROM_MEM[11227] = 8'h05;
ROM_MEM[11228] = 8'h05;
ROM_MEM[11229] = 8'h01;
ROM_MEM[11230] = 8'hB1;
ROM_MEM[11231] = 8'h06;
ROM_MEM[11232] = 8'h07;
ROM_MEM[11233] = 8'h01;
ROM_MEM[11234] = 8'hCF;
ROM_MEM[11235] = 8'h07;
ROM_MEM[11236] = 8'h03;
ROM_MEM[11237] = 8'h01;
ROM_MEM[11238] = 8'h3C;
ROM_MEM[11239] = 8'h01;
ROM_MEM[11240] = 8'h0A;
ROM_MEM[11241] = 8'h01;
ROM_MEM[11242] = 8'h40;
ROM_MEM[11243] = 8'h02;
ROM_MEM[11244] = 8'h0D;
ROM_MEM[11245] = 8'h01;
ROM_MEM[11246] = 8'h55;
ROM_MEM[11247] = 8'h03;
ROM_MEM[11248] = 8'h09;
ROM_MEM[11249] = 8'h01;
ROM_MEM[11250] = 8'h7D;
ROM_MEM[11251] = 8'h04;
ROM_MEM[11252] = 8'h08;
ROM_MEM[11253] = 8'h01;
ROM_MEM[11254] = 8'hA2;
ROM_MEM[11255] = 8'h05;
ROM_MEM[11256] = 8'h06;
ROM_MEM[11257] = 8'h01;
ROM_MEM[11258] = 8'hCB;
ROM_MEM[11259] = 8'h06;
ROM_MEM[11260] = 8'h03;
ROM_MEM[11261] = 8'h01;
ROM_MEM[11262] = 8'hF1;
ROM_MEM[11263] = 8'h07;
ROM_MEM[11264] = 8'h03;
ROM_MEM[11265] = 8'h06;
ROM_MEM[11266] = 8'hAF;
ROM_MEM[11267] = 8'hFF;
ROM_MEM[11268] = 8'h03;
ROM_MEM[11269] = 8'h06;
ROM_MEM[11270] = 8'hAB;
ROM_MEM[11271] = 8'hFE;
ROM_MEM[11272] = 8'h02;
ROM_MEM[11273] = 8'h08;
ROM_MEM[11274] = 8'hA4;
ROM_MEM[11275] = 8'hFD;
ROM_MEM[11276] = 8'h00;
ROM_MEM[11277] = 8'hC0;
ROM_MEM[11278] = 8'h01;
ROM_MEM[11279] = 8'hEC;
ROM_MEM[11280] = 8'hFF;
ROM_MEM[11281] = 8'h24;
ROM_MEM[11282] = 8'h02;
ROM_MEM[11283] = 8'h2C;
ROM_MEM[11284] = 8'hFF;
ROM_MEM[11285] = 8'h06;
ROM_MEM[11286] = 8'h02;
ROM_MEM[11287] = 8'h0A;
ROM_MEM[11288] = 8'h01;
ROM_MEM[11289] = 8'h03;
ROM_MEM[11290] = 8'h04;
ROM_MEM[11291] = 8'h0F;
ROM_MEM[11292] = 8'h01;
ROM_MEM[11293] = 8'h02;
ROM_MEM[11294] = 8'h06;
ROM_MEM[11295] = 8'h12;
ROM_MEM[11296] = 8'hFF;
ROM_MEM[11297] = 8'h02;
ROM_MEM[11298] = 8'h08;
ROM_MEM[11299] = 8'h10;
ROM_MEM[11300] = 8'hFF;
ROM_MEM[11301] = 8'h02;
ROM_MEM[11302] = 8'h0A;
ROM_MEM[11303] = 8'h0E;
ROM_MEM[11304] = 8'hFF;
ROM_MEM[11305] = 8'h01;
ROM_MEM[11306] = 8'h0E;
ROM_MEM[11307] = 8'h0C;
ROM_MEM[11308] = 8'h00;
ROM_MEM[11309] = 8'h01;
ROM_MEM[11310] = 8'hBC;
ROM_MEM[11311] = 8'h82;
ROM_MEM[11312] = 8'h00;
ROM_MEM[11313] = 8'h01;
ROM_MEM[11314] = 8'h08;
ROM_MEM[11315] = 8'h83;
ROM_MEM[11316] = 8'h00;
ROM_MEM[11317] = 8'h01;
ROM_MEM[11318] = 8'h08;
ROM_MEM[11319] = 8'h84;
ROM_MEM[11320] = 8'h00;
ROM_MEM[11321] = 8'h04;
ROM_MEM[11322] = 8'h08;
ROM_MEM[11323] = 8'h85;
ROM_MEM[11324] = 8'h01;
ROM_MEM[11325] = 8'h02;
ROM_MEM[11326] = 8'h06;
ROM_MEM[11327] = 8'h89;
ROM_MEM[11328] = 8'h01;
ROM_MEM[11329] = 8'h02;
ROM_MEM[11330] = 8'h04;
ROM_MEM[11331] = 8'h8B;
ROM_MEM[11332] = 8'h01;
ROM_MEM[11333] = 8'h01;
ROM_MEM[11334] = 8'h06;
ROM_MEM[11335] = 8'h8D;
ROM_MEM[11336] = 8'h00;
ROM_MEM[11337] = 8'h02;
ROM_MEM[11338] = 8'h04;
ROM_MEM[11339] = 8'h8E;
ROM_MEM[11340] = 8'h01;
ROM_MEM[11341] = 8'h07;
ROM_MEM[11342] = 8'h02;
ROM_MEM[11343] = 8'h8E;
ROM_MEM[11344] = 8'hFF;
ROM_MEM[11345] = 8'h02;
ROM_MEM[11346] = 8'h04;
ROM_MEM[11347] = 8'h87;
ROM_MEM[11348] = 8'hFF;
ROM_MEM[11349] = 8'h01;
ROM_MEM[11350] = 8'h06;
ROM_MEM[11351] = 8'h85;
ROM_MEM[11352] = 8'h00;
ROM_MEM[11353] = 8'h01;
ROM_MEM[11354] = 8'h04;
ROM_MEM[11355] = 8'h84;
ROM_MEM[11356] = 8'h00;
ROM_MEM[11357] = 8'h01;
ROM_MEM[11358] = 8'h06;
ROM_MEM[11359] = 8'h83;
ROM_MEM[11360] = 8'h00;
ROM_MEM[11361] = 8'h01;
ROM_MEM[11362] = 8'h10;
ROM_MEM[11363] = 8'h82;
ROM_MEM[11364] = 8'h00;
ROM_MEM[11365] = 8'h01;
ROM_MEM[11366] = 8'h1A;
ROM_MEM[11367] = 8'h81;
ROM_MEM[11368] = 8'h00;
ROM_MEM[11369] = 8'h00;
ROM_MEM[11370] = 8'hA0;
ROM_MEM[11371] = 8'h01;
ROM_MEM[11372] = 8'hE5;
ROM_MEM[11373] = 8'hFF;
ROM_MEM[11374] = 8'h30;
ROM_MEM[11375] = 8'h02;
ROM_MEM[11376] = 8'h45;
ROM_MEM[11377] = 8'hFF;
ROM_MEM[11378] = 8'h0E;
ROM_MEM[11379] = 8'h02;
ROM_MEM[11380] = 8'h16;
ROM_MEM[11381] = 8'h01;
ROM_MEM[11382] = 8'h01;
ROM_MEM[11383] = 8'h42;
ROM_MEM[11384] = 8'h16;
ROM_MEM[11385] = 8'h00;
ROM_MEM[11386] = 8'h01;
ROM_MEM[11387] = 8'hA0;
ROM_MEM[11388] = 8'hC1;
ROM_MEM[11389] = 8'h00;
ROM_MEM[11390] = 8'h07;
ROM_MEM[11391] = 8'h08;
ROM_MEM[11392] = 8'hC1;
ROM_MEM[11393] = 8'h01;
ROM_MEM[11394] = 8'h02;
ROM_MEM[11395] = 8'h06;
ROM_MEM[11396] = 8'hC9;
ROM_MEM[11397] = 8'h01;
ROM_MEM[11398] = 8'h02;
ROM_MEM[11399] = 8'h04;
ROM_MEM[11400] = 8'hCB;
ROM_MEM[11401] = 8'h01;
ROM_MEM[11402] = 8'h01;
ROM_MEM[11403] = 8'h06;
ROM_MEM[11404] = 8'hCD;
ROM_MEM[11405] = 8'h00;
ROM_MEM[11406] = 8'h02;
ROM_MEM[11407] = 8'h04;
ROM_MEM[11408] = 8'hCE;
ROM_MEM[11409] = 8'h01;
ROM_MEM[11410] = 8'h0E;
ROM_MEM[11411] = 8'h02;
ROM_MEM[11412] = 8'hCE;
ROM_MEM[11413] = 8'hFF;
ROM_MEM[11414] = 8'h01;
ROM_MEM[11415] = 8'h42;
ROM_MEM[11416] = 8'hC0;
ROM_MEM[11417] = 8'h00;
ROM_MEM[11418] = 8'h00;
ROM_MEM[11419] = 8'h1E;
ROM_MEM[11420] = 8'h01;
ROM_MEM[11421] = 8'h51;
ROM_MEM[11422] = 8'hFE;
ROM_MEM[11423] = 8'h1E;
ROM_MEM[11424] = 8'h01;
ROM_MEM[11425] = 8'hA2;
ROM_MEM[11426] = 8'h02;
ROM_MEM[11427] = 8'h01;
ROM_MEM[11428] = 8'h1E;
ROM_MEM[11429] = 8'hAA;
ROM_MEM[11430] = 8'h00;
ROM_MEM[11431] = 8'h00;
ROM_MEM[11432] = 8'h08;
ROM_MEM[11433] = 8'h32;
ROM_MEM[11434] = 8'h66;
ROM_MEM[11435] = 8'h00;
ROM_MEM[11436] = 8'h01;
ROM_MEM[11437] = 8'h28;
ROM_MEM[11438] = 8'hAA;
ROM_MEM[11439] = 8'h00;
ROM_MEM[11440] = 8'h00;
ROM_MEM[11441] = 8'h08;
ROM_MEM[11442] = 8'h32;
ROM_MEM[11443] = 8'h5B;
ROM_MEM[11444] = 8'h00;
ROM_MEM[11445] = 8'h02;
ROM_MEM[11446] = 8'h28;
ROM_MEM[11447] = 8'hA0;
ROM_MEM[11448] = 8'h0A;
ROM_MEM[11449] = 8'h00;
ROM_MEM[11450] = 8'h08;
ROM_MEM[11451] = 8'h32;
ROM_MEM[11452] = 8'h51;
ROM_MEM[11453] = 8'h00;
ROM_MEM[11454] = 8'h01;
ROM_MEM[11455] = 8'h50;
ROM_MEM[11456] = 8'hA0;
ROM_MEM[11457] = 8'h00;
ROM_MEM[11458] = 8'h01;
ROM_MEM[11459] = 8'h28;
ROM_MEM[11460] = 8'hAA;
ROM_MEM[11461] = 8'h00;
ROM_MEM[11462] = 8'h00;
ROM_MEM[11463] = 8'h08;
ROM_MEM[11464] = 8'h32;
ROM_MEM[11465] = 8'h48;
ROM_MEM[11466] = 8'h00;
ROM_MEM[11467] = 8'h01;
ROM_MEM[11468] = 8'h78;
ROM_MEM[11469] = 8'hA0;
ROM_MEM[11470] = 8'h00;
ROM_MEM[11471] = 8'h01;
ROM_MEM[11472] = 8'h28;
ROM_MEM[11473] = 8'hAA;
ROM_MEM[11474] = 8'h00;
ROM_MEM[11475] = 8'h00;
ROM_MEM[11476] = 8'h01;
ROM_MEM[11477] = 8'hA0;
ROM_MEM[11478] = 8'hA0;
ROM_MEM[11479] = 8'h00;
ROM_MEM[11480] = 8'h02;
ROM_MEM[11481] = 8'h0F;
ROM_MEM[11482] = 8'hAA;
ROM_MEM[11483] = 8'hF6;
ROM_MEM[11484] = 8'h02;
ROM_MEM[11485] = 8'h0F;
ROM_MEM[11486] = 8'hAA;
ROM_MEM[11487] = 8'hF6;
ROM_MEM[11488] = 8'h00;
ROM_MEM[11489] = 8'h01;
ROM_MEM[11490] = 8'hDC;
ROM_MEM[11491] = 8'hA0;
ROM_MEM[11492] = 8'h00;
ROM_MEM[11493] = 8'h02;
ROM_MEM[11494] = 8'h0F;
ROM_MEM[11495] = 8'hAA;
ROM_MEM[11496] = 8'hF6;
ROM_MEM[11497] = 8'h02;
ROM_MEM[11498] = 8'h0F;
ROM_MEM[11499] = 8'hAA;
ROM_MEM[11500] = 8'hF6;
ROM_MEM[11501] = 8'h00;
ROM_MEM[11502] = 8'h02;
ROM_MEM[11503] = 8'h8C;
ROM_MEM[11504] = 8'hA0;
ROM_MEM[11505] = 8'h00;
ROM_MEM[11506] = 8'h02;
ROM_MEM[11507] = 8'h0F;
ROM_MEM[11508] = 8'hAA;
ROM_MEM[11509] = 8'hF6;
ROM_MEM[11510] = 8'h02;
ROM_MEM[11511] = 8'h0F;
ROM_MEM[11512] = 8'hAA;
ROM_MEM[11513] = 8'hF6;
ROM_MEM[11514] = 8'h00;
ROM_MEM[11515] = 8'h02;
ROM_MEM[11516] = 8'hAA;
ROM_MEM[11517] = 8'hA0;
ROM_MEM[11518] = 8'h00;
ROM_MEM[11519] = 8'h02;
ROM_MEM[11520] = 8'h0F;
ROM_MEM[11521] = 8'hAA;
ROM_MEM[11522] = 8'hF6;
ROM_MEM[11523] = 8'h02;
ROM_MEM[11524] = 8'h0F;
ROM_MEM[11525] = 8'hAA;
ROM_MEM[11526] = 8'hF6;
ROM_MEM[11527] = 8'h00;
ROM_MEM[11528] = 8'h01;
ROM_MEM[11529] = 8'hF0;
ROM_MEM[11530] = 8'h0C;
ROM_MEM[11531] = 8'h00;
ROM_MEM[11532] = 8'h01;
ROM_MEM[11533] = 8'h09;
ROM_MEM[11534] = 8'h0C;
ROM_MEM[11535] = 8'h00;
ROM_MEM[11536] = 8'h01;
ROM_MEM[11537] = 8'h2A;
ROM_MEM[11538] = 8'h0F;
ROM_MEM[11539] = 8'h00;
ROM_MEM[11540] = 8'h01;
ROM_MEM[11541] = 8'h05;
ROM_MEM[11542] = 8'h0C;
ROM_MEM[11543] = 8'h00;
ROM_MEM[11544] = 8'h01;
ROM_MEM[11545] = 8'h15;
ROM_MEM[11546] = 8'h14;
ROM_MEM[11547] = 8'h00;
ROM_MEM[11548] = 8'h01;
ROM_MEM[11549] = 8'h0C;
ROM_MEM[11550] = 8'h0C;
ROM_MEM[11551] = 8'h00;
ROM_MEM[11552] = 8'h01;
ROM_MEM[11553] = 8'h11;
ROM_MEM[11554] = 8'h0F;
ROM_MEM[11555] = 8'h00;
ROM_MEM[11556] = 8'h01;
ROM_MEM[11557] = 8'h0D;
ROM_MEM[11558] = 8'h0C;
ROM_MEM[11559] = 8'h00;
ROM_MEM[11560] = 8'h01;
ROM_MEM[11561] = 8'h15;
ROM_MEM[11562] = 8'h14;
ROM_MEM[11563] = 8'h00;
ROM_MEM[11564] = 8'h01;
ROM_MEM[11565] = 8'h0C;
ROM_MEM[11566] = 8'h0C;
ROM_MEM[11567] = 8'h00;
ROM_MEM[11568] = 8'h01;
ROM_MEM[11569] = 8'h22;
ROM_MEM[11570] = 8'h0F;
ROM_MEM[11571] = 8'h00;
ROM_MEM[11572] = 8'h01;
ROM_MEM[11573] = 8'h0D;
ROM_MEM[11574] = 8'h17;
ROM_MEM[11575] = 8'h00;
ROM_MEM[11576] = 8'h01;
ROM_MEM[11577] = 8'h07;
ROM_MEM[11578] = 8'h15;
ROM_MEM[11579] = 8'h00;
ROM_MEM[11580] = 8'h02;
ROM_MEM[11581] = 8'h01;
ROM_MEM[11582] = 8'h14;
ROM_MEM[11583] = 8'hFF;
ROM_MEM[11584] = 8'h01;
ROM_MEM[11585] = 8'h03;
ROM_MEM[11586] = 8'h15;
ROM_MEM[11587] = 8'h00;
ROM_MEM[11588] = 8'h02;
ROM_MEM[11589] = 8'h01;
ROM_MEM[11590] = 8'h13;
ROM_MEM[11591] = 8'hFF;
ROM_MEM[11592] = 8'h02;
ROM_MEM[11593] = 8'h01;
ROM_MEM[11594] = 8'h10;
ROM_MEM[11595] = 8'hFE;
ROM_MEM[11596] = 8'h02;
ROM_MEM[11597] = 8'h01;
ROM_MEM[11598] = 8'h0D;
ROM_MEM[11599] = 8'hFF;
ROM_MEM[11600] = 8'h01;
ROM_MEM[11601] = 8'h02;
ROM_MEM[11602] = 8'h0B;
ROM_MEM[11603] = 8'h00;
ROM_MEM[11604] = 8'h03;
ROM_MEM[11605] = 8'h01;
ROM_MEM[11606] = 8'h09;
ROM_MEM[11607] = 8'hFF;
ROM_MEM[11608] = 8'h01;
ROM_MEM[11609] = 8'h0E;
ROM_MEM[11610] = 8'h06;
ROM_MEM[11611] = 8'h00;
ROM_MEM[11612] = 8'h01;
ROM_MEM[11613] = 8'h01;
ROM_MEM[11614] = 8'h07;
ROM_MEM[11615] = 8'h00;
ROM_MEM[11616] = 8'h01;
ROM_MEM[11617] = 8'h02;
ROM_MEM[11618] = 8'h08;
ROM_MEM[11619] = 8'h00;
ROM_MEM[11620] = 8'h06;
ROM_MEM[11621] = 8'h01;
ROM_MEM[11622] = 8'h09;
ROM_MEM[11623] = 8'h01;
ROM_MEM[11624] = 8'h01;
ROM_MEM[11625] = 8'h02;
ROM_MEM[11626] = 8'h10;
ROM_MEM[11627] = 8'h00;
ROM_MEM[11628] = 8'h01;
ROM_MEM[11629] = 8'h01;
ROM_MEM[11630] = 8'h12;
ROM_MEM[11631] = 8'h00;
ROM_MEM[11632] = 8'h01;
ROM_MEM[11633] = 8'hF0;
ROM_MEM[11634] = 8'hA0;
ROM_MEM[11635] = 8'h00;
ROM_MEM[11636] = 8'h01;
ROM_MEM[11637] = 8'h05;
ROM_MEM[11638] = 8'hAA;
ROM_MEM[11639] = 8'h00;
ROM_MEM[11640] = 8'h01;
ROM_MEM[11641] = 8'h04;
ROM_MEM[11642] = 8'h00;
ROM_MEM[11643] = 8'h00;
ROM_MEM[11644] = 8'h01;
ROM_MEM[11645] = 8'h0A;
ROM_MEM[11646] = 8'hAB;
ROM_MEM[11647] = 8'h00;
ROM_MEM[11648] = 8'h01;
ROM_MEM[11649] = 8'h20;
ROM_MEM[11650] = 8'h00;
ROM_MEM[11651] = 8'h00;
ROM_MEM[11652] = 8'h01;
ROM_MEM[11653] = 8'h05;
ROM_MEM[11654] = 8'hAB;
ROM_MEM[11655] = 8'h00;
ROM_MEM[11656] = 8'h01;
ROM_MEM[11657] = 8'h0A;
ROM_MEM[11658] = 8'hAC;
ROM_MEM[11659] = 8'h00;
ROM_MEM[11660] = 8'h01;
ROM_MEM[11661] = 8'h0B;
ROM_MEM[11662] = 8'h00;
ROM_MEM[11663] = 8'h00;
ROM_MEM[11664] = 8'h01;
ROM_MEM[11665] = 8'h06;
ROM_MEM[11666] = 8'hAB;
ROM_MEM[11667] = 8'h00;
ROM_MEM[11668] = 8'h01;
ROM_MEM[11669] = 8'h06;
ROM_MEM[11670] = 8'h00;
ROM_MEM[11671] = 8'h00;
ROM_MEM[11672] = 8'h01;
ROM_MEM[11673] = 8'h09;
ROM_MEM[11674] = 8'hAC;
ROM_MEM[11675] = 8'h00;
ROM_MEM[11676] = 8'h01;
ROM_MEM[11677] = 8'h08;
ROM_MEM[11678] = 8'h00;
ROM_MEM[11679] = 8'h00;
ROM_MEM[11680] = 8'h01;
ROM_MEM[11681] = 8'h08;
ROM_MEM[11682] = 8'hAA;
ROM_MEM[11683] = 8'h00;
ROM_MEM[11684] = 8'h01;
ROM_MEM[11685] = 8'h05;
ROM_MEM[11686] = 8'h00;
ROM_MEM[11687] = 8'h00;
ROM_MEM[11688] = 8'h01;
ROM_MEM[11689] = 8'h0A;
ROM_MEM[11690] = 8'hAC;
ROM_MEM[11691] = 8'h00;
ROM_MEM[11692] = 8'h01;
ROM_MEM[11693] = 8'h0B;
ROM_MEM[11694] = 8'h00;
ROM_MEM[11695] = 8'h00;
ROM_MEM[11696] = 8'h01;
ROM_MEM[11697] = 8'h06;
ROM_MEM[11698] = 8'hAB;
ROM_MEM[11699] = 8'h00;
ROM_MEM[11700] = 8'h01;
ROM_MEM[11701] = 8'h06;
ROM_MEM[11702] = 8'h00;
ROM_MEM[11703] = 8'h00;
ROM_MEM[11704] = 8'h01;
ROM_MEM[11705] = 8'h09;
ROM_MEM[11706] = 8'hAC;
ROM_MEM[11707] = 8'h00;
ROM_MEM[11708] = 8'h01;
ROM_MEM[11709] = 8'h19;
ROM_MEM[11710] = 8'h00;
ROM_MEM[11711] = 8'h00;
ROM_MEM[11712] = 8'h03;
ROM_MEM[11713] = 8'h01;
ROM_MEM[11714] = 8'hA2;
ROM_MEM[11715] = 8'h01;
ROM_MEM[11716] = 8'h04;
ROM_MEM[11717] = 8'h01;
ROM_MEM[11718] = 8'hA6;
ROM_MEM[11719] = 8'h01;
ROM_MEM[11720] = 8'h03;
ROM_MEM[11721] = 8'h01;
ROM_MEM[11722] = 8'hA8;
ROM_MEM[11723] = 8'hFF;
ROM_MEM[11724] = 8'h01;
ROM_MEM[11725] = 8'h02;
ROM_MEM[11726] = 8'hA5;
ROM_MEM[11727] = 8'h00;
ROM_MEM[11728] = 8'h02;
ROM_MEM[11729] = 8'h01;
ROM_MEM[11730] = 8'hA7;
ROM_MEM[11731] = 8'h03;
ROM_MEM[11732] = 8'h01;
ROM_MEM[11733] = 8'h04;
ROM_MEM[11734] = 8'hAC;
ROM_MEM[11735] = 8'h00;
ROM_MEM[11736] = 8'h03;
ROM_MEM[11737] = 8'h01;
ROM_MEM[11738] = 8'hAB;
ROM_MEM[11739] = 8'hFD;
ROM_MEM[11740] = 8'h02;
ROM_MEM[11741] = 8'h02;
ROM_MEM[11742] = 8'hA3;
ROM_MEM[11743] = 8'hFF;
ROM_MEM[11744] = 8'h02;
ROM_MEM[11745] = 8'h01;
ROM_MEM[11746] = 8'hA3;
ROM_MEM[11747] = 8'h06;
ROM_MEM[11748] = 8'h01;
ROM_MEM[11749] = 8'h06;
ROM_MEM[11750] = 8'hAD;
ROM_MEM[11751] = 8'h00;
ROM_MEM[11752] = 8'h01;
ROM_MEM[11753] = 8'h01;
ROM_MEM[11754] = 8'hAC;
ROM_MEM[11755] = 8'h00;
ROM_MEM[11756] = 8'h01;
ROM_MEM[11757] = 8'h02;
ROM_MEM[11758] = 8'hAA;
ROM_MEM[11759] = 8'h00;
ROM_MEM[11760] = 8'h01;
ROM_MEM[11761] = 8'h01;
ROM_MEM[11762] = 8'hA9;
ROM_MEM[11763] = 8'h00;
ROM_MEM[11764] = 8'h01;
ROM_MEM[11765] = 8'h08;
ROM_MEM[11766] = 8'hA8;
ROM_MEM[11767] = 8'h00;
ROM_MEM[11768] = 8'h01;
ROM_MEM[11769] = 8'h06;
ROM_MEM[11770] = 8'hA7;
ROM_MEM[11771] = 8'h00;
ROM_MEM[11772] = 8'h01;
ROM_MEM[11773] = 8'h05;
ROM_MEM[11774] = 8'hA8;
ROM_MEM[11775] = 8'h00;
ROM_MEM[11776] = 8'h01;
ROM_MEM[11777] = 8'h02;
ROM_MEM[11778] = 8'hA9;
ROM_MEM[11779] = 8'h00;
ROM_MEM[11780] = 8'h01;
ROM_MEM[11781] = 8'h01;
ROM_MEM[11782] = 8'hA8;
ROM_MEM[11783] = 8'h00;
ROM_MEM[11784] = 8'h03;
ROM_MEM[11785] = 8'h01;
ROM_MEM[11786] = 8'hA6;
ROM_MEM[11787] = 8'hFF;
ROM_MEM[11788] = 8'h00;
ROM_MEM[11789] = 8'h01;
ROM_MEM[11790] = 8'hC0;
ROM_MEM[11791] = 8'h12;
ROM_MEM[11792] = 8'h00;
ROM_MEM[11793] = 8'h01;
ROM_MEM[11794] = 8'h01;
ROM_MEM[11795] = 8'h12;
ROM_MEM[11796] = 8'h00;
ROM_MEM[11797] = 8'h01;
ROM_MEM[11798] = 8'h06;
ROM_MEM[11799] = 8'h13;
ROM_MEM[11800] = 8'h00;
ROM_MEM[11801] = 8'h01;
ROM_MEM[11802] = 8'h0A;
ROM_MEM[11803] = 8'h14;
ROM_MEM[11804] = 8'h00;
ROM_MEM[11805] = 8'h01;
ROM_MEM[11806] = 8'h18;
ROM_MEM[11807] = 8'h0B;
ROM_MEM[11808] = 8'h00;
ROM_MEM[11809] = 8'h01;
ROM_MEM[11810] = 8'h0E;
ROM_MEM[11811] = 8'h18;
ROM_MEM[11812] = 8'h00;
ROM_MEM[11813] = 8'h01;
ROM_MEM[11814] = 8'h04;
ROM_MEM[11815] = 8'h15;
ROM_MEM[11816] = 8'h00;
ROM_MEM[11817] = 8'h01;
ROM_MEM[11818] = 8'h04;
ROM_MEM[11819] = 8'h0F;
ROM_MEM[11820] = 8'h00;
ROM_MEM[11821] = 8'h01;
ROM_MEM[11822] = 8'h05;
ROM_MEM[11823] = 8'h0B;
ROM_MEM[11824] = 8'h00;
ROM_MEM[11825] = 8'h01;
ROM_MEM[11826] = 8'h0A;
ROM_MEM[11827] = 8'h05;
ROM_MEM[11828] = 8'h00;
ROM_MEM[11829] = 8'h02;
ROM_MEM[11830] = 8'h01;
ROM_MEM[11831] = 8'h0E;
ROM_MEM[11832] = 8'h03;
ROM_MEM[11833] = 8'h06;
ROM_MEM[11834] = 8'h01;
ROM_MEM[11835] = 8'h13;
ROM_MEM[11836] = 8'h01;
ROM_MEM[11837] = 8'h01;
ROM_MEM[11838] = 8'h01;
ROM_MEM[11839] = 8'h17;
ROM_MEM[11840] = 8'h00;
ROM_MEM[11841] = 8'h01;
ROM_MEM[11842] = 8'h02;
ROM_MEM[11843] = 8'h18;
ROM_MEM[11844] = 8'h00;
ROM_MEM[11845] = 8'h01;
ROM_MEM[11846] = 8'h20;
ROM_MEM[11847] = 8'h16;
ROM_MEM[11848] = 8'h00;
ROM_MEM[11849] = 8'h02;
ROM_MEM[11850] = 8'h01;
ROM_MEM[11851] = 8'h3F;
ROM_MEM[11852] = 8'hFA;
ROM_MEM[11853] = 8'h03;
ROM_MEM[11854] = 8'h01;
ROM_MEM[11855] = 8'h36;
ROM_MEM[11856] = 8'hFE;
ROM_MEM[11857] = 8'h02;
ROM_MEM[11858] = 8'h01;
ROM_MEM[11859] = 8'h2F;
ROM_MEM[11860] = 8'hFC;
ROM_MEM[11861] = 8'h02;
ROM_MEM[11862] = 8'h01;
ROM_MEM[11863] = 8'h29;
ROM_MEM[11864] = 8'hFF;
ROM_MEM[11865] = 8'h03;
ROM_MEM[11866] = 8'h01;
ROM_MEM[11867] = 8'h26;
ROM_MEM[11868] = 8'hFF;
ROM_MEM[11869] = 8'h01;
ROM_MEM[11870] = 8'h01;
ROM_MEM[11871] = 8'h22;
ROM_MEM[11872] = 8'h00;
ROM_MEM[11873] = 8'h03;
ROM_MEM[11874] = 8'h01;
ROM_MEM[11875] = 8'h22;
ROM_MEM[11876] = 8'hFE;
ROM_MEM[11877] = 8'h05;
ROM_MEM[11878] = 8'h01;
ROM_MEM[11879] = 8'h1D;
ROM_MEM[11880] = 8'hFF;
ROM_MEM[11881] = 8'h01;
ROM_MEM[11882] = 8'h04;
ROM_MEM[11883] = 8'h18;
ROM_MEM[11884] = 8'h00;
ROM_MEM[11885] = 8'h01;
ROM_MEM[11886] = 8'h02;
ROM_MEM[11887] = 8'h17;
ROM_MEM[11888] = 8'h00;
ROM_MEM[11889] = 8'h01;
ROM_MEM[11890] = 8'h01;
ROM_MEM[11891] = 8'h16;
ROM_MEM[11892] = 8'h00;
ROM_MEM[11893] = 8'h01;
ROM_MEM[11894] = 8'h04;
ROM_MEM[11895] = 8'h15;
ROM_MEM[11896] = 8'h00;
ROM_MEM[11897] = 8'h01;
ROM_MEM[11898] = 8'h01;
ROM_MEM[11899] = 8'h14;
ROM_MEM[11900] = 8'h00;
ROM_MEM[11901] = 8'h02;
ROM_MEM[11902] = 8'h03;
ROM_MEM[11903] = 8'h13;
ROM_MEM[11904] = 8'hFF;
ROM_MEM[11905] = 8'h01;
ROM_MEM[11906] = 8'h02;
ROM_MEM[11907] = 8'h11;
ROM_MEM[11908] = 8'h00;
ROM_MEM[11909] = 8'h02;
ROM_MEM[11910] = 8'h01;
ROM_MEM[11911] = 8'h10;
ROM_MEM[11912] = 8'h01;
ROM_MEM[11913] = 8'h01;
ROM_MEM[11914] = 8'h06;
ROM_MEM[11915] = 8'h10;
ROM_MEM[11916] = 8'h00;
ROM_MEM[11917] = 8'h01;
ROM_MEM[11918] = 8'h04;
ROM_MEM[11919] = 8'h0F;
ROM_MEM[11920] = 8'h00;
ROM_MEM[11921] = 8'h01;
ROM_MEM[11922] = 8'h15;
ROM_MEM[11923] = 8'h0E;
ROM_MEM[11924] = 8'h00;
ROM_MEM[11925] = 8'h01;
ROM_MEM[11926] = 8'h0E;
ROM_MEM[11927] = 8'h13;
ROM_MEM[11928] = 8'h00;
ROM_MEM[11929] = 8'h01;
ROM_MEM[11930] = 8'h03;
ROM_MEM[11931] = 8'h0B;
ROM_MEM[11932] = 8'h00;
ROM_MEM[11933] = 8'h01;
ROM_MEM[11934] = 8'h0D;
ROM_MEM[11935] = 8'h10;
ROM_MEM[11936] = 8'h00;
ROM_MEM[11937] = 8'h01;
ROM_MEM[11938] = 8'h05;
ROM_MEM[11939] = 8'h10;
ROM_MEM[11940] = 8'h00;
ROM_MEM[11941] = 8'h01;
ROM_MEM[11942] = 8'h0E;
ROM_MEM[11943] = 8'h09;
ROM_MEM[11944] = 8'h00;
ROM_MEM[11945] = 8'h01;
ROM_MEM[11946] = 8'h0C;
ROM_MEM[11947] = 8'h13;
ROM_MEM[11948] = 8'h00;
ROM_MEM[11949] = 8'h01;
ROM_MEM[11950] = 8'hC0;
ROM_MEM[11951] = 8'hA0;
ROM_MEM[11952] = 8'h00;
ROM_MEM[11953] = 8'h01;
ROM_MEM[11954] = 8'h01;
ROM_MEM[11955] = 8'hA8;
ROM_MEM[11956] = 8'h00;
ROM_MEM[11957] = 8'h01;
ROM_MEM[11958] = 8'h07;
ROM_MEM[11959] = 8'hAA;
ROM_MEM[11960] = 8'h00;
ROM_MEM[11961] = 8'h01;
ROM_MEM[11962] = 8'h09;
ROM_MEM[11963] = 8'hA0;
ROM_MEM[11964] = 8'h00;
ROM_MEM[11965] = 8'h02;
ROM_MEM[11966] = 8'h0C;
ROM_MEM[11967] = 8'hA8;
ROM_MEM[11968] = 8'hF8;
ROM_MEM[11969] = 8'h01;
ROM_MEM[11970] = 8'h06;
ROM_MEM[11971] = 8'hAD;
ROM_MEM[11972] = 8'h00;
ROM_MEM[11973] = 8'h01;
ROM_MEM[11974] = 8'h03;
ROM_MEM[11975] = 8'hA0;
ROM_MEM[11976] = 8'h00;
ROM_MEM[11977] = 8'h01;
ROM_MEM[11978] = 8'h05;
ROM_MEM[11979] = 8'hAD;
ROM_MEM[11980] = 8'h00;
ROM_MEM[11981] = 8'h01;
ROM_MEM[11982] = 8'h01;
ROM_MEM[11983] = 8'hAA;
ROM_MEM[11984] = 8'h00;
ROM_MEM[11985] = 8'h01;
ROM_MEM[11986] = 8'h03;
ROM_MEM[11987] = 8'hA0;
ROM_MEM[11988] = 8'h00;
ROM_MEM[11989] = 8'h01;
ROM_MEM[11990] = 8'h04;
ROM_MEM[11991] = 8'hAA;
ROM_MEM[11992] = 8'h00;
ROM_MEM[11993] = 8'h01;
ROM_MEM[11994] = 8'h01;
ROM_MEM[11995] = 8'hA9;
ROM_MEM[11996] = 8'h00;
ROM_MEM[11997] = 8'h01;
ROM_MEM[11998] = 8'h0E;
ROM_MEM[11999] = 8'hA0;
ROM_MEM[12000] = 8'h00;
ROM_MEM[12001] = 8'h03;
ROM_MEM[12002] = 8'h01;
ROM_MEM[12003] = 8'hAA;
ROM_MEM[12004] = 8'h01;
ROM_MEM[12005] = 8'h01;
ROM_MEM[12006] = 8'h06;
ROM_MEM[12007] = 8'hAD;
ROM_MEM[12008] = 8'h00;
ROM_MEM[12009] = 8'h01;
ROM_MEM[12010] = 8'h02;
ROM_MEM[12011] = 8'hAC;
ROM_MEM[12012] = 8'h00;
ROM_MEM[12013] = 8'h01;
ROM_MEM[12014] = 8'h01;
ROM_MEM[12015] = 8'hA5;
ROM_MEM[12016] = 8'h00;
ROM_MEM[12017] = 8'h01;
ROM_MEM[12018] = 8'h1F;
ROM_MEM[12019] = 8'hA0;
ROM_MEM[12020] = 8'h00;
ROM_MEM[12021] = 8'h01;
ROM_MEM[12022] = 8'h01;
ROM_MEM[12023] = 8'hA6;
ROM_MEM[12024] = 8'h00;
ROM_MEM[12025] = 8'h01;
ROM_MEM[12026] = 8'h02;
ROM_MEM[12027] = 8'hA7;
ROM_MEM[12028] = 8'h00;
ROM_MEM[12029] = 8'h01;
ROM_MEM[12030] = 8'h04;
ROM_MEM[12031] = 8'hA8;
ROM_MEM[12032] = 8'h00;
ROM_MEM[12033] = 8'h01;
ROM_MEM[12034] = 8'h05;
ROM_MEM[12035] = 8'hA9;
ROM_MEM[12036] = 8'h00;
ROM_MEM[12037] = 8'h01;
ROM_MEM[12038] = 8'h02;
ROM_MEM[12039] = 8'hAA;
ROM_MEM[12040] = 8'h00;
ROM_MEM[12041] = 8'h02;
ROM_MEM[12042] = 8'h01;
ROM_MEM[12043] = 8'hAB;
ROM_MEM[12044] = 8'h01;
ROM_MEM[12045] = 8'h01;
ROM_MEM[12046] = 8'h01;
ROM_MEM[12047] = 8'hAB;
ROM_MEM[12048] = 8'h00;
ROM_MEM[12049] = 8'h01;
ROM_MEM[12050] = 8'h02;
ROM_MEM[12051] = 8'hAC;
ROM_MEM[12052] = 8'h00;
ROM_MEM[12053] = 8'h02;
ROM_MEM[12054] = 8'h01;
ROM_MEM[12055] = 8'hAB;
ROM_MEM[12056] = 8'hFF;
ROM_MEM[12057] = 8'h01;
ROM_MEM[12058] = 8'h20;
ROM_MEM[12059] = 8'hA9;
ROM_MEM[12060] = 8'h00;
ROM_MEM[12061] = 8'h01;
ROM_MEM[12062] = 8'h0C;
ROM_MEM[12063] = 8'hA8;
ROM_MEM[12064] = 8'h00;
ROM_MEM[12065] = 8'h01;
ROM_MEM[12066] = 8'h09;
ROM_MEM[12067] = 8'hA0;
ROM_MEM[12068] = 8'h00;
ROM_MEM[12069] = 8'h01;
ROM_MEM[12070] = 8'h0E;
ROM_MEM[12071] = 8'hAA;
ROM_MEM[12072] = 8'h00;
ROM_MEM[12073] = 8'h01;
ROM_MEM[12074] = 8'h03;
ROM_MEM[12075] = 8'hA9;
ROM_MEM[12076] = 8'h00;
ROM_MEM[12077] = 8'h01;
ROM_MEM[12078] = 8'h0D;
ROM_MEM[12079] = 8'hAA;
ROM_MEM[12080] = 8'h00;
ROM_MEM[12081] = 8'h01;
ROM_MEM[12082] = 8'h05;
ROM_MEM[12083] = 8'hA0;
ROM_MEM[12084] = 8'h00;
ROM_MEM[12085] = 8'h01;
ROM_MEM[12086] = 8'h1A;
ROM_MEM[12087] = 8'hA6;
ROM_MEM[12088] = 8'h00;
ROM_MEM[12089] = 8'h00;
ROM_MEM[12090] = 8'h02;
ROM_MEM[12091] = 8'h01;
ROM_MEM[12092] = 8'h3B;
ROM_MEM[12093] = 8'hD8;
ROM_MEM[12094] = 8'h01;
ROM_MEM[12095] = 8'h01;
ROM_MEM[12096] = 8'h0D;
ROM_MEM[12097] = 8'h00;
ROM_MEM[12098] = 8'h03;
ROM_MEM[12099] = 8'h01;
ROM_MEM[12100] = 8'h07;
ROM_MEM[12101] = 8'hFE;
ROM_MEM[12102] = 8'h01;
ROM_MEM[12103] = 8'h07;
ROM_MEM[12104] = 8'h04;
ROM_MEM[12105] = 8'h00;
ROM_MEM[12106] = 8'h02;
ROM_MEM[12107] = 8'h02;
ROM_MEM[12108] = 8'h05;
ROM_MEM[12109] = 8'h01;
ROM_MEM[12110] = 8'h01;
ROM_MEM[12111] = 8'h01;
ROM_MEM[12112] = 8'h08;
ROM_MEM[12113] = 8'h00;
ROM_MEM[12114] = 8'h01;
ROM_MEM[12115] = 8'h03;
ROM_MEM[12116] = 8'h0A;
ROM_MEM[12117] = 8'h00;
ROM_MEM[12118] = 8'h02;
ROM_MEM[12119] = 8'h01;
ROM_MEM[12120] = 8'h0C;
ROM_MEM[12121] = 8'h01;
ROM_MEM[12122] = 8'h01;
ROM_MEM[12123] = 8'h02;
ROM_MEM[12124] = 8'h0E;
ROM_MEM[12125] = 8'h00;
ROM_MEM[12126] = 8'h01;
ROM_MEM[12127] = 8'h04;
ROM_MEM[12128] = 8'h0D;
ROM_MEM[12129] = 8'h00;
ROM_MEM[12130] = 8'h02;
ROM_MEM[12131] = 8'h02;
ROM_MEM[12132] = 8'h0E;
ROM_MEM[12133] = 8'hFF;
ROM_MEM[12134] = 8'h01;
ROM_MEM[12135] = 8'h01;
ROM_MEM[12136] = 8'h0C;
ROM_MEM[12137] = 8'h00;
ROM_MEM[12138] = 8'h01;
ROM_MEM[12139] = 8'h03;
ROM_MEM[12140] = 8'h0D;
ROM_MEM[12141] = 8'h00;
ROM_MEM[12142] = 8'h01;
ROM_MEM[12143] = 8'h01;
ROM_MEM[12144] = 8'h70;
ROM_MEM[12145] = 8'h00;
ROM_MEM[12146] = 8'h01;
ROM_MEM[12147] = 8'h07;
ROM_MEM[12148] = 8'h10;
ROM_MEM[12149] = 8'h00;
ROM_MEM[12150] = 8'h03;
ROM_MEM[12151] = 8'h01;
ROM_MEM[12152] = 8'h09;
ROM_MEM[12153] = 8'hFE;
ROM_MEM[12154] = 8'h02;
ROM_MEM[12155] = 8'h01;
ROM_MEM[12156] = 8'h04;
ROM_MEM[12157] = 8'hFF;
ROM_MEM[12158] = 8'h02;
ROM_MEM[12159] = 8'h01;
ROM_MEM[12160] = 8'h03;
ROM_MEM[12161] = 8'h02;
ROM_MEM[12162] = 8'h01;
ROM_MEM[12163] = 8'h02;
ROM_MEM[12164] = 8'h07;
ROM_MEM[12165] = 8'h00;
ROM_MEM[12166] = 8'h01;
ROM_MEM[12167] = 8'h09;
ROM_MEM[12168] = 8'h03;
ROM_MEM[12169] = 8'h00;
ROM_MEM[12170] = 8'h01;
ROM_MEM[12171] = 8'h03;
ROM_MEM[12172] = 8'h07;
ROM_MEM[12173] = 8'h00;
ROM_MEM[12174] = 8'h02;
ROM_MEM[12175] = 8'h01;
ROM_MEM[12176] = 8'h05;
ROM_MEM[12177] = 8'h03;
ROM_MEM[12178] = 8'h02;
ROM_MEM[12179] = 8'h01;
ROM_MEM[12180] = 8'h0C;
ROM_MEM[12181] = 8'h05;
ROM_MEM[12182] = 8'h02;
ROM_MEM[12183] = 8'h01;
ROM_MEM[12184] = 8'h18;
ROM_MEM[12185] = 8'hFD;
ROM_MEM[12186] = 8'h01;
ROM_MEM[12187] = 8'h02;
ROM_MEM[12188] = 8'h0A;
ROM_MEM[12189] = 8'h00;
ROM_MEM[12190] = 8'h02;
ROM_MEM[12191] = 8'h01;
ROM_MEM[12192] = 8'h10;
ROM_MEM[12193] = 8'h02;
ROM_MEM[12194] = 8'h01;
ROM_MEM[12195] = 8'h02;
ROM_MEM[12196] = 8'h1D;
ROM_MEM[12197] = 8'h00;
ROM_MEM[12198] = 8'h02;
ROM_MEM[12199] = 8'h01;
ROM_MEM[12200] = 8'h25;
ROM_MEM[12201] = 8'hFC;
ROM_MEM[12202] = 8'h02;
ROM_MEM[12203] = 8'h01;
ROM_MEM[12204] = 8'h19;
ROM_MEM[12205] = 8'hF7;
ROM_MEM[12206] = 8'h01;
ROM_MEM[12207] = 8'h01;
ROM_MEM[12208] = 8'h0C;
ROM_MEM[12209] = 8'h00;
ROM_MEM[12210] = 8'h01;
ROM_MEM[12211] = 8'h04;
ROM_MEM[12212] = 8'h0A;
ROM_MEM[12213] = 8'h00;
ROM_MEM[12214] = 8'h01;
ROM_MEM[12215] = 8'h05;
ROM_MEM[12216] = 8'h09;
ROM_MEM[12217] = 8'h00;
ROM_MEM[12218] = 8'h01;
ROM_MEM[12219] = 8'h01;
ROM_MEM[12220] = 8'h0B;
ROM_MEM[12221] = 8'h00;
ROM_MEM[12222] = 8'h01;
ROM_MEM[12223] = 8'h02;
ROM_MEM[12224] = 8'h0C;
ROM_MEM[12225] = 8'h00;
ROM_MEM[12226] = 8'h02;
ROM_MEM[12227] = 8'h01;
ROM_MEM[12228] = 8'h0B;
ROM_MEM[12229] = 8'hFE;
ROM_MEM[12230] = 8'h02;
ROM_MEM[12231] = 8'h01;
ROM_MEM[12232] = 8'h08;
ROM_MEM[12233] = 8'h08;
ROM_MEM[12234] = 8'h02;
ROM_MEM[12235] = 8'h01;
ROM_MEM[12236] = 8'h2A;
ROM_MEM[12237] = 8'h03;
ROM_MEM[12238] = 8'h01;
ROM_MEM[12239] = 8'h01;
ROM_MEM[12240] = 8'h29;
ROM_MEM[12241] = 8'h00;
ROM_MEM[12242] = 8'h01;
ROM_MEM[12243] = 8'h05;
ROM_MEM[12244] = 8'h28;
ROM_MEM[12245] = 8'h00;
ROM_MEM[12246] = 8'h02;
ROM_MEM[12247] = 8'h01;
ROM_MEM[12248] = 8'h26;
ROM_MEM[12249] = 8'h1A;
ROM_MEM[12250] = 8'h01;
ROM_MEM[12251] = 8'h01;
ROM_MEM[12252] = 8'h1B;
ROM_MEM[12253] = 8'h00;
ROM_MEM[12254] = 8'h03;
ROM_MEM[12255] = 8'h01;
ROM_MEM[12256] = 8'h0D;
ROM_MEM[12257] = 8'hFF;
ROM_MEM[12258] = 8'h01;
ROM_MEM[12259] = 8'h06;
ROM_MEM[12260] = 8'h0A;
ROM_MEM[12261] = 8'h00;
ROM_MEM[12262] = 8'h01;
ROM_MEM[12263] = 8'h03;
ROM_MEM[12264] = 8'h0B;
ROM_MEM[12265] = 8'h00;
ROM_MEM[12266] = 8'h02;
ROM_MEM[12267] = 8'h01;
ROM_MEM[12268] = 8'h0C;
ROM_MEM[12269] = 8'h01;
ROM_MEM[12270] = 8'h01;
ROM_MEM[12271] = 8'h05;
ROM_MEM[12272] = 8'h0E;
ROM_MEM[12273] = 8'h00;
ROM_MEM[12274] = 8'h03;
ROM_MEM[12275] = 8'h01;
ROM_MEM[12276] = 8'h0F;
ROM_MEM[12277] = 8'hFF;
ROM_MEM[12278] = 8'h01;
ROM_MEM[12279] = 8'h02;
ROM_MEM[12280] = 8'h0B;
ROM_MEM[12281] = 8'h00;
ROM_MEM[12282] = 8'h02;
ROM_MEM[12283] = 8'h05;
ROM_MEM[12284] = 8'h09;
ROM_MEM[12285] = 8'hFF;
ROM_MEM[12286] = 8'h02;
ROM_MEM[12287] = 8'h01;
ROM_MEM[12288] = 8'h0A;
ROM_MEM[12289] = 8'h01;
ROM_MEM[12290] = 8'h02;
ROM_MEM[12291] = 8'h01;
ROM_MEM[12292] = 8'h0E;
ROM_MEM[12293] = 8'h02;
ROM_MEM[12294] = 8'h01;
ROM_MEM[12295] = 8'h01;
ROM_MEM[12296] = 8'h16;
ROM_MEM[12297] = 8'h00;
ROM_MEM[12298] = 8'h02;
ROM_MEM[12299] = 8'h02;
ROM_MEM[12300] = 8'h19;
ROM_MEM[12301] = 8'hF1;
ROM_MEM[12302] = 8'h02;
ROM_MEM[12303] = 8'h01;
ROM_MEM[12304] = 8'h0D;
ROM_MEM[12305] = 8'hFC;
ROM_MEM[12306] = 8'h02;
ROM_MEM[12307] = 8'h01;
ROM_MEM[12308] = 8'h0C;
ROM_MEM[12309] = 8'h01;
ROM_MEM[12310] = 8'h01;
ROM_MEM[12311] = 8'h01;
ROM_MEM[12312] = 8'h11;
ROM_MEM[12313] = 8'h00;
ROM_MEM[12314] = 8'h01;
ROM_MEM[12315] = 8'h02;
ROM_MEM[12316] = 8'h12;
ROM_MEM[12317] = 8'h00;
ROM_MEM[12318] = 8'h02;
ROM_MEM[12319] = 8'h01;
ROM_MEM[12320] = 8'hA1;
ROM_MEM[12321] = 8'h01;
ROM_MEM[12322] = 8'h04;
ROM_MEM[12323] = 8'h01;
ROM_MEM[12324] = 8'hA5;
ROM_MEM[12325] = 8'hFF;
ROM_MEM[12326] = 8'h03;
ROM_MEM[12327] = 8'h01;
ROM_MEM[12328] = 8'hA1;
ROM_MEM[12329] = 8'h01;
ROM_MEM[12330] = 8'h01;
ROM_MEM[12331] = 8'h03;
ROM_MEM[12332] = 8'hA3;
ROM_MEM[12333] = 8'h00;
ROM_MEM[12334] = 8'h02;
ROM_MEM[12335] = 8'h01;
ROM_MEM[12336] = 8'hA4;
ROM_MEM[12337] = 8'h01;
ROM_MEM[12338] = 8'h01;
ROM_MEM[12339] = 8'h01;
ROM_MEM[12340] = 8'hA7;
ROM_MEM[12341] = 8'h00;
ROM_MEM[12342] = 8'h01;
ROM_MEM[12343] = 8'h0B;
ROM_MEM[12344] = 8'hAA;
ROM_MEM[12345] = 8'h00;
ROM_MEM[12346] = 8'h02;
ROM_MEM[12347] = 8'h01;
ROM_MEM[12348] = 8'hA7;
ROM_MEM[12349] = 8'hFA;
ROM_MEM[12350] = 8'h01;
ROM_MEM[12351] = 8'h0A;
ROM_MEM[12352] = 8'hA1;
ROM_MEM[12353] = 8'h00;
ROM_MEM[12354] = 8'h01;
ROM_MEM[12355] = 8'h06;
ROM_MEM[12356] = 8'hA0;
ROM_MEM[12357] = 8'h00;
ROM_MEM[12358] = 8'h01;
ROM_MEM[12359] = 8'h01;
ROM_MEM[12360] = 8'hA8;
ROM_MEM[12361] = 8'h00;
ROM_MEM[12362] = 8'h01;
ROM_MEM[12363] = 8'h02;
ROM_MEM[12364] = 8'hAA;
ROM_MEM[12365] = 8'h00;
ROM_MEM[12366] = 8'h02;
ROM_MEM[12367] = 8'h01;
ROM_MEM[12368] = 8'hA7;
ROM_MEM[12369] = 8'hFB;
ROM_MEM[12370] = 8'h01;
ROM_MEM[12371] = 8'h05;
ROM_MEM[12372] = 8'hA1;
ROM_MEM[12373] = 8'h00;
ROM_MEM[12374] = 8'h02;
ROM_MEM[12375] = 8'h02;
ROM_MEM[12376] = 8'hA0;
ROM_MEM[12377] = 8'h01;
ROM_MEM[12378] = 8'h01;
ROM_MEM[12379] = 8'h03;
ROM_MEM[12380] = 8'hA1;
ROM_MEM[12381] = 8'h00;
ROM_MEM[12382] = 8'h02;
ROM_MEM[12383] = 8'h02;
ROM_MEM[12384] = 8'hA1;
ROM_MEM[12385] = 8'hFF;
ROM_MEM[12386] = 8'h02;
ROM_MEM[12387] = 8'h01;
ROM_MEM[12388] = 8'hA1;
ROM_MEM[12389] = 8'h03;
ROM_MEM[12390] = 8'h01;
ROM_MEM[12391] = 8'h05;
ROM_MEM[12392] = 8'hAA;
ROM_MEM[12393] = 8'h00;
ROM_MEM[12394] = 8'h02;
ROM_MEM[12395] = 8'h01;
ROM_MEM[12396] = 8'hA5;
ROM_MEM[12397] = 8'hFC;
ROM_MEM[12398] = 8'h01;
ROM_MEM[12399] = 8'h02;
ROM_MEM[12400] = 8'hA1;
ROM_MEM[12401] = 8'h00;
ROM_MEM[12402] = 8'h02;
ROM_MEM[12403] = 8'h01;
ROM_MEM[12404] = 8'hA0;
ROM_MEM[12405] = 8'h05;
ROM_MEM[12406] = 8'h01;
ROM_MEM[12407] = 8'h06;
ROM_MEM[12408] = 8'hAA;
ROM_MEM[12409] = 8'h00;
ROM_MEM[12410] = 8'h02;
ROM_MEM[12411] = 8'h01;
ROM_MEM[12412] = 8'hA7;
ROM_MEM[12413] = 8'hFF;
ROM_MEM[12414] = 8'h02;
ROM_MEM[12415] = 8'h01;
ROM_MEM[12416] = 8'hA7;
ROM_MEM[12417] = 8'h02;
ROM_MEM[12418] = 8'h01;
ROM_MEM[12419] = 8'h05;
ROM_MEM[12420] = 8'hAA;
ROM_MEM[12421] = 8'h00;
ROM_MEM[12422] = 8'h02;
ROM_MEM[12423] = 8'h01;
ROM_MEM[12424] = 8'hA9;
ROM_MEM[12425] = 8'hF9;
ROM_MEM[12426] = 8'h01;
ROM_MEM[12427] = 8'h03;
ROM_MEM[12428] = 8'hA1;
ROM_MEM[12429] = 8'h00;
ROM_MEM[12430] = 8'h03;
ROM_MEM[12431] = 8'h01;
ROM_MEM[12432] = 8'hA2;
ROM_MEM[12433] = 8'h03;
ROM_MEM[12434] = 8'h01;
ROM_MEM[12435] = 8'h04;
ROM_MEM[12436] = 8'hAA;
ROM_MEM[12437] = 8'h00;
ROM_MEM[12438] = 8'h03;
ROM_MEM[12439] = 8'h01;
ROM_MEM[12440] = 8'hA8;
ROM_MEM[12441] = 8'hFD;
ROM_MEM[12442] = 8'h01;
ROM_MEM[12443] = 8'h01;
ROM_MEM[12444] = 8'hA1;
ROM_MEM[12445] = 8'h00;
ROM_MEM[12446] = 8'h01;
ROM_MEM[12447] = 8'h06;
ROM_MEM[12448] = 8'hAA;
ROM_MEM[12449] = 8'h00;
ROM_MEM[12450] = 8'h01;
ROM_MEM[12451] = 8'h02;
ROM_MEM[12452] = 8'hA7;
ROM_MEM[12453] = 8'h00;
ROM_MEM[12454] = 8'h02;
ROM_MEM[12455] = 8'h01;
ROM_MEM[12456] = 8'hA5;
ROM_MEM[12457] = 8'hFD;
ROM_MEM[12458] = 8'h01;
ROM_MEM[12459] = 8'h02;
ROM_MEM[12460] = 8'hA1;
ROM_MEM[12461] = 8'h00;
ROM_MEM[12462] = 8'h02;
ROM_MEM[12463] = 8'h01;
ROM_MEM[12464] = 8'hA1;
ROM_MEM[12465] = 8'h08;
ROM_MEM[12466] = 8'h01;
ROM_MEM[12467] = 8'h05;
ROM_MEM[12468] = 8'hAA;
ROM_MEM[12469] = 8'h00;
ROM_MEM[12470] = 8'h02;
ROM_MEM[12471] = 8'h01;
ROM_MEM[12472] = 8'hA4;
ROM_MEM[12473] = 8'hFD;
ROM_MEM[12474] = 8'h02;
ROM_MEM[12475] = 8'h01;
ROM_MEM[12476] = 8'hA1;
ROM_MEM[12477] = 8'h01;
ROM_MEM[12478] = 8'h02;
ROM_MEM[12479] = 8'h01;
ROM_MEM[12480] = 8'hA4;
ROM_MEM[12481] = 8'h04;
ROM_MEM[12482] = 8'h01;
ROM_MEM[12483] = 8'h03;
ROM_MEM[12484] = 8'hAA;
ROM_MEM[12485] = 8'h00;
ROM_MEM[12486] = 8'h01;
ROM_MEM[12487] = 8'h01;
ROM_MEM[12488] = 8'hA9;
ROM_MEM[12489] = 8'h00;
ROM_MEM[12490] = 8'h01;
ROM_MEM[12491] = 8'h03;
ROM_MEM[12492] = 8'hA7;
ROM_MEM[12493] = 8'h00;
ROM_MEM[12494] = 8'h01;
ROM_MEM[12495] = 8'h01;
ROM_MEM[12496] = 8'hA9;
ROM_MEM[12497] = 8'h00;
ROM_MEM[12498] = 8'h01;
ROM_MEM[12499] = 8'h07;
ROM_MEM[12500] = 8'hAA;
ROM_MEM[12501] = 8'h00;
ROM_MEM[12502] = 8'h02;
ROM_MEM[12503] = 8'h01;
ROM_MEM[12504] = 8'hA8;
ROM_MEM[12505] = 8'hFD;
ROM_MEM[12506] = 8'h01;
ROM_MEM[12507] = 8'h09;
ROM_MEM[12508] = 8'hA1;
ROM_MEM[12509] = 8'h00;
ROM_MEM[12510] = 8'h00;
ROM_MEM[12511] = 8'h01;
ROM_MEM[12512] = 8'h06;
ROM_MEM[12513] = 8'h08;
ROM_MEM[12514] = 8'h00;
ROM_MEM[12515] = 8'h01;
ROM_MEM[12516] = 8'h04;
ROM_MEM[12517] = 8'h09;
ROM_MEM[12518] = 8'h00;
ROM_MEM[12519] = 8'h01;
ROM_MEM[12520] = 8'h02;
ROM_MEM[12521] = 8'h08;
ROM_MEM[12522] = 8'h00;
ROM_MEM[12523] = 8'h01;
ROM_MEM[12524] = 8'h01;
ROM_MEM[12525] = 8'h09;
ROM_MEM[12526] = 8'h00;
ROM_MEM[12527] = 8'h01;
ROM_MEM[12528] = 8'h03;
ROM_MEM[12529] = 8'h0A;
ROM_MEM[12530] = 8'h00;
ROM_MEM[12531] = 8'h01;
ROM_MEM[12532] = 8'h01;
ROM_MEM[12533] = 8'h0B;
ROM_MEM[12534] = 8'h00;
ROM_MEM[12535] = 8'h01;
ROM_MEM[12536] = 8'h02;
ROM_MEM[12537] = 8'h0A;
ROM_MEM[12538] = 8'h00;
ROM_MEM[12539] = 8'h01;
ROM_MEM[12540] = 8'h01;
ROM_MEM[12541] = 8'h0B;
ROM_MEM[12542] = 8'h00;
ROM_MEM[12543] = 8'h01;
ROM_MEM[12544] = 8'h03;
ROM_MEM[12545] = 8'h0A;
ROM_MEM[12546] = 8'h00;
ROM_MEM[12547] = 8'h01;
ROM_MEM[12548] = 8'h01;
ROM_MEM[12549] = 8'h0B;
ROM_MEM[12550] = 8'h00;
ROM_MEM[12551] = 8'h02;
ROM_MEM[12552] = 8'h02;
ROM_MEM[12553] = 8'h0C;
ROM_MEM[12554] = 8'hFF;
ROM_MEM[12555] = 8'h01;
ROM_MEM[12556] = 8'h03;
ROM_MEM[12557] = 8'h0A;
ROM_MEM[12558] = 8'h00;
ROM_MEM[12559] = 8'h01;
ROM_MEM[12560] = 8'h05;
ROM_MEM[12561] = 8'h0B;
ROM_MEM[12562] = 8'h00;
ROM_MEM[12563] = 8'h01;
ROM_MEM[12564] = 8'h14;
ROM_MEM[12565] = 8'h0A;
ROM_MEM[12566] = 8'h00;
ROM_MEM[12567] = 8'h01;
ROM_MEM[12568] = 8'h02;
ROM_MEM[12569] = 8'h0B;
ROM_MEM[12570] = 8'h00;
ROM_MEM[12571] = 8'h01;
ROM_MEM[12572] = 8'h01;
ROM_MEM[12573] = 8'h0D;
ROM_MEM[12574] = 8'h00;
ROM_MEM[12575] = 8'h01;
ROM_MEM[12576] = 8'h02;
ROM_MEM[12577] = 8'h0C;
ROM_MEM[12578] = 8'h00;
ROM_MEM[12579] = 8'h01;
ROM_MEM[12580] = 8'h04;
ROM_MEM[12581] = 8'h0D;
ROM_MEM[12582] = 8'h00;
ROM_MEM[12583] = 8'h01;
ROM_MEM[12584] = 8'h01;
ROM_MEM[12585] = 8'h0E;
ROM_MEM[12586] = 8'h00;
ROM_MEM[12587] = 8'h01;
ROM_MEM[12588] = 8'h02;
ROM_MEM[12589] = 8'h0F;
ROM_MEM[12590] = 8'h00;
ROM_MEM[12591] = 8'h02;
ROM_MEM[12592] = 8'h01;
ROM_MEM[12593] = 8'h10;
ROM_MEM[12594] = 8'h01;
ROM_MEM[12595] = 8'h01;
ROM_MEM[12596] = 8'h02;
ROM_MEM[12597] = 8'h12;
ROM_MEM[12598] = 8'h00;
ROM_MEM[12599] = 8'h01;
ROM_MEM[12600] = 8'h01;
ROM_MEM[12601] = 8'h14;
ROM_MEM[12602] = 8'h00;
ROM_MEM[12603] = 8'h01;
ROM_MEM[12604] = 8'h05;
ROM_MEM[12605] = 8'h13;
ROM_MEM[12606] = 8'h00;
ROM_MEM[12607] = 8'h01;
ROM_MEM[12608] = 8'h02;
ROM_MEM[12609] = 8'h14;
ROM_MEM[12610] = 8'h00;
ROM_MEM[12611] = 8'h01;
ROM_MEM[12612] = 8'h04;
ROM_MEM[12613] = 8'h13;
ROM_MEM[12614] = 8'h00;
ROM_MEM[12615] = 8'h01;
ROM_MEM[12616] = 8'h02;
ROM_MEM[12617] = 8'h14;
ROM_MEM[12618] = 8'h00;
ROM_MEM[12619] = 8'h01;
ROM_MEM[12620] = 8'h01;
ROM_MEM[12621] = 8'h13;
ROM_MEM[12622] = 8'h00;
ROM_MEM[12623] = 8'h01;
ROM_MEM[12624] = 8'h04;
ROM_MEM[12625] = 8'h12;
ROM_MEM[12626] = 8'h00;
ROM_MEM[12627] = 8'h01;
ROM_MEM[12628] = 8'h03;
ROM_MEM[12629] = 8'h11;
ROM_MEM[12630] = 8'h00;
ROM_MEM[12631] = 8'h01;
ROM_MEM[12632] = 8'h02;
ROM_MEM[12633] = 8'h10;
ROM_MEM[12634] = 8'h00;
ROM_MEM[12635] = 8'h01;
ROM_MEM[12636] = 8'h09;
ROM_MEM[12637] = 8'h0F;
ROM_MEM[12638] = 8'h00;
ROM_MEM[12639] = 8'h01;
ROM_MEM[12640] = 8'h04;
ROM_MEM[12641] = 8'h10;
ROM_MEM[12642] = 8'h00;
ROM_MEM[12643] = 8'h01;
ROM_MEM[12644] = 8'h03;
ROM_MEM[12645] = 8'h11;
ROM_MEM[12646] = 8'h00;
ROM_MEM[12647] = 8'h01;
ROM_MEM[12648] = 8'h05;
ROM_MEM[12649] = 8'h12;
ROM_MEM[12650] = 8'h00;
ROM_MEM[12651] = 8'h01;
ROM_MEM[12652] = 8'h01;
ROM_MEM[12653] = 8'h13;
ROM_MEM[12654] = 8'h00;
ROM_MEM[12655] = 8'h01;
ROM_MEM[12656] = 8'h02;
ROM_MEM[12657] = 8'h23;
ROM_MEM[12658] = 8'hFF;
ROM_MEM[12659] = 8'h01;
ROM_MEM[12660] = 8'h04;
ROM_MEM[12661] = 8'h21;
ROM_MEM[12662] = 8'h00;
ROM_MEM[12663] = 8'h01;
ROM_MEM[12664] = 8'h03;
ROM_MEM[12665] = 8'h23;
ROM_MEM[12666] = 8'h00;
ROM_MEM[12667] = 8'h01;
ROM_MEM[12668] = 8'h02;
ROM_MEM[12669] = 8'h24;
ROM_MEM[12670] = 8'h00;
ROM_MEM[12671] = 8'h02;
ROM_MEM[12672] = 8'h01;
ROM_MEM[12673] = 8'h25;
ROM_MEM[12674] = 8'h01;
ROM_MEM[12675] = 8'h01;
ROM_MEM[12676] = 8'h02;
ROM_MEM[12677] = 8'h27;
ROM_MEM[12678] = 8'h00;
ROM_MEM[12679] = 8'h01;
ROM_MEM[12680] = 8'h01;
ROM_MEM[12681] = 8'h26;
ROM_MEM[12682] = 8'h00;
ROM_MEM[12683] = 8'h01;
ROM_MEM[12684] = 8'h03;
ROM_MEM[12685] = 8'h25;
ROM_MEM[12686] = 8'h00;
ROM_MEM[12687] = 8'h01;
ROM_MEM[12688] = 8'h02;
ROM_MEM[12689] = 8'h24;
ROM_MEM[12690] = 8'h00;
ROM_MEM[12691] = 8'h01;
ROM_MEM[12692] = 8'h06;
ROM_MEM[12693] = 8'h23;
ROM_MEM[12694] = 8'h00;
ROM_MEM[12695] = 8'h02;
ROM_MEM[12696] = 8'h01;
ROM_MEM[12697] = 8'h22;
ROM_MEM[12698] = 8'hFF;
ROM_MEM[12699] = 8'h02;
ROM_MEM[12700] = 8'h01;
ROM_MEM[12701] = 8'h23;
ROM_MEM[12702] = 8'hFF;
ROM_MEM[12703] = 8'h01;
ROM_MEM[12704] = 8'h03;
ROM_MEM[12705] = 8'h21;
ROM_MEM[12706] = 8'h00;
ROM_MEM[12707] = 8'h02;
ROM_MEM[12708] = 8'h02;
ROM_MEM[12709] = 8'h22;
ROM_MEM[12710] = 8'hFF;
ROM_MEM[12711] = 8'h01;
ROM_MEM[12712] = 8'h01;
ROM_MEM[12713] = 8'h22;
ROM_MEM[12714] = 8'h00;
ROM_MEM[12715] = 8'h01;
ROM_MEM[12716] = 8'h02;
ROM_MEM[12717] = 8'h23;
ROM_MEM[12718] = 8'h00;
ROM_MEM[12719] = 8'h03;
ROM_MEM[12720] = 8'h01;
ROM_MEM[12721] = 8'h24;
ROM_MEM[12722] = 8'h01;
ROM_MEM[12723] = 8'h01;
ROM_MEM[12724] = 8'h04;
ROM_MEM[12725] = 8'h27;
ROM_MEM[12726] = 8'h00;
ROM_MEM[12727] = 8'h02;
ROM_MEM[12728] = 8'h01;
ROM_MEM[12729] = 8'h29;
ROM_MEM[12730] = 8'h02;
ROM_MEM[12731] = 8'h01;
ROM_MEM[12732] = 8'h02;
ROM_MEM[12733] = 8'h2E;
ROM_MEM[12734] = 8'h00;
ROM_MEM[12735] = 8'h01;
ROM_MEM[12736] = 8'h01;
ROM_MEM[12737] = 8'h31;
ROM_MEM[12738] = 8'h00;
ROM_MEM[12739] = 8'h01;
ROM_MEM[12740] = 8'h02;
ROM_MEM[12741] = 8'h2F;
ROM_MEM[12742] = 8'h00;
ROM_MEM[12743] = 8'h02;
ROM_MEM[12744] = 8'h01;
ROM_MEM[12745] = 8'h33;
ROM_MEM[12746] = 8'h06;
ROM_MEM[12747] = 8'h02;
ROM_MEM[12748] = 8'h01;
ROM_MEM[12749] = 8'h36;
ROM_MEM[12750] = 8'hFC;
ROM_MEM[12751] = 8'h02;
ROM_MEM[12752] = 8'h01;
ROM_MEM[12753] = 8'h2C;
ROM_MEM[12754] = 8'h06;
ROM_MEM[12755] = 8'h02;
ROM_MEM[12756] = 8'h01;
ROM_MEM[12757] = 8'h31;
ROM_MEM[12758] = 8'h01;
ROM_MEM[12759] = 8'h02;
ROM_MEM[12760] = 8'h01;
ROM_MEM[12761] = 8'h30;
ROM_MEM[12762] = 8'h02;
ROM_MEM[12763] = 8'h02;
ROM_MEM[12764] = 8'h01;
ROM_MEM[12765] = 8'h30;
ROM_MEM[12766] = 8'h01;
ROM_MEM[12767] = 8'h01;
ROM_MEM[12768] = 8'h02;
ROM_MEM[12769] = 8'h32;
ROM_MEM[12770] = 8'h00;
ROM_MEM[12771] = 8'h01;
ROM_MEM[12772] = 8'h01;
ROM_MEM[12773] = 8'h33;
ROM_MEM[12774] = 8'h00;
ROM_MEM[12775] = 8'h01;
ROM_MEM[12776] = 8'h03;
ROM_MEM[12777] = 8'h34;
ROM_MEM[12778] = 8'h00;
ROM_MEM[12779] = 8'h01;
ROM_MEM[12780] = 8'h02;
ROM_MEM[12781] = 8'h36;
ROM_MEM[12782] = 8'h00;
ROM_MEM[12783] = 8'h01;
ROM_MEM[12784] = 8'h01;
ROM_MEM[12785] = 8'h38;
ROM_MEM[12786] = 8'h00;
ROM_MEM[12787] = 8'h01;
ROM_MEM[12788] = 8'h03;
ROM_MEM[12789] = 8'h37;
ROM_MEM[12790] = 8'h00;
ROM_MEM[12791] = 8'h02;
ROM_MEM[12792] = 8'h01;
ROM_MEM[12793] = 8'h38;
ROM_MEM[12794] = 8'hFC;
ROM_MEM[12795] = 8'h01;
ROM_MEM[12796] = 8'h01;
ROM_MEM[12797] = 8'h35;
ROM_MEM[12798] = 8'h00;
ROM_MEM[12799] = 8'h01;
ROM_MEM[12800] = 8'h02;
ROM_MEM[12801] = 8'h40;
ROM_MEM[12802] = 8'h00;
ROM_MEM[12803] = 8'h02;
ROM_MEM[12804] = 8'h01;
ROM_MEM[12805] = 8'h45;
ROM_MEM[12806] = 8'hFD;
ROM_MEM[12807] = 8'h03;
ROM_MEM[12808] = 8'h01;
ROM_MEM[12809] = 8'h35;
ROM_MEM[12810] = 8'h08;
ROM_MEM[12811] = 8'h02;
ROM_MEM[12812] = 8'h01;
ROM_MEM[12813] = 8'h46;
ROM_MEM[12814] = 8'hFE;
ROM_MEM[12815] = 8'h02;
ROM_MEM[12816] = 8'h01;
ROM_MEM[12817] = 8'h40;
ROM_MEM[12818] = 8'h02;
ROM_MEM[12819] = 8'h01;
ROM_MEM[12820] = 8'h04;
ROM_MEM[12821] = 8'h43;
ROM_MEM[12822] = 8'h00;
ROM_MEM[12823] = 8'h02;
ROM_MEM[12824] = 8'h01;
ROM_MEM[12825] = 8'h42;
ROM_MEM[12826] = 8'hFE;
ROM_MEM[12827] = 8'h02;
ROM_MEM[12828] = 8'h01;
ROM_MEM[12829] = 8'h36;
ROM_MEM[12830] = 8'hFB;
ROM_MEM[12831] = 8'h01;
ROM_MEM[12832] = 8'h1D;
ROM_MEM[12833] = 8'hA1;
ROM_MEM[12834] = 8'h00;
ROM_MEM[12835] = 8'h01;
ROM_MEM[12836] = 8'h05;
ROM_MEM[12837] = 8'hA2;
ROM_MEM[12838] = 8'h00;
ROM_MEM[12839] = 8'h01;
ROM_MEM[12840] = 8'h14;
ROM_MEM[12841] = 8'hA1;
ROM_MEM[12842] = 8'h00;
ROM_MEM[12843] = 8'h01;
ROM_MEM[12844] = 8'h02;
ROM_MEM[12845] = 8'hA2;
ROM_MEM[12846] = 8'h00;
ROM_MEM[12847] = 8'h01;
ROM_MEM[12848] = 8'h03;
ROM_MEM[12849] = 8'hA3;
ROM_MEM[12850] = 8'h00;
ROM_MEM[12851] = 8'h01;
ROM_MEM[12852] = 8'h03;
ROM_MEM[12853] = 8'hA7;
ROM_MEM[12854] = 8'h00;
ROM_MEM[12855] = 8'h02;
ROM_MEM[12856] = 8'h02;
ROM_MEM[12857] = 8'hA8;
ROM_MEM[12858] = 8'h01;
ROM_MEM[12859] = 8'h01;
ROM_MEM[12860] = 8'h01;
ROM_MEM[12861] = 8'hA8;
ROM_MEM[12862] = 8'h00;
ROM_MEM[12863] = 8'h01;
ROM_MEM[12864] = 8'h02;
ROM_MEM[12865] = 8'hA9;
ROM_MEM[12866] = 8'h00;
ROM_MEM[12867] = 8'h02;
ROM_MEM[12868] = 8'h01;
ROM_MEM[12869] = 8'hA8;
ROM_MEM[12870] = 8'h01;
ROM_MEM[12871] = 8'h01;
ROM_MEM[12872] = 8'h0F;
ROM_MEM[12873] = 8'hAA;
ROM_MEM[12874] = 8'h00;
ROM_MEM[12875] = 8'h02;
ROM_MEM[12876] = 8'h01;
ROM_MEM[12877] = 8'hA9;
ROM_MEM[12878] = 8'hFF;
ROM_MEM[12879] = 8'h02;
ROM_MEM[12880] = 8'h01;
ROM_MEM[12881] = 8'hA6;
ROM_MEM[12882] = 8'hFE;
ROM_MEM[12883] = 8'h01;
ROM_MEM[12884] = 8'h07;
ROM_MEM[12885] = 8'hA3;
ROM_MEM[12886] = 8'h00;
ROM_MEM[12887] = 8'h01;
ROM_MEM[12888] = 8'h01;
ROM_MEM[12889] = 8'hA2;
ROM_MEM[12890] = 8'h00;
ROM_MEM[12891] = 8'h01;
ROM_MEM[12892] = 8'h14;
ROM_MEM[12893] = 8'hA1;
ROM_MEM[12894] = 8'h00;
ROM_MEM[12895] = 8'h01;
ROM_MEM[12896] = 8'h1A;
ROM_MEM[12897] = 8'hAA;
ROM_MEM[12898] = 8'h00;
ROM_MEM[12899] = 8'h01;
ROM_MEM[12900] = 8'h0E;
ROM_MEM[12901] = 8'hA8;
ROM_MEM[12902] = 8'h00;
ROM_MEM[12903] = 8'h01;
ROM_MEM[12904] = 8'h05;
ROM_MEM[12905] = 8'hAA;
ROM_MEM[12906] = 8'h00;
ROM_MEM[12907] = 8'h03;
ROM_MEM[12908] = 8'h01;
ROM_MEM[12909] = 8'hA8;
ROM_MEM[12910] = 8'hFF;
ROM_MEM[12911] = 8'h02;
ROM_MEM[12912] = 8'h01;
ROM_MEM[12913] = 8'hA4;
ROM_MEM[12914] = 8'hFD;
ROM_MEM[12915] = 8'h02;
ROM_MEM[12916] = 8'h04;
ROM_MEM[12917] = 8'hA1;
ROM_MEM[12918] = 8'h01;
ROM_MEM[12919] = 8'h01;
ROM_MEM[12920] = 8'h01;
ROM_MEM[12921] = 8'hA2;
ROM_MEM[12922] = 8'h00;
ROM_MEM[12923] = 8'h01;
ROM_MEM[12924] = 8'h0B;
ROM_MEM[12925] = 8'hA1;
ROM_MEM[12926] = 8'h00;
ROM_MEM[12927] = 8'h03;
ROM_MEM[12928] = 8'h02;
ROM_MEM[12929] = 8'hA2;
ROM_MEM[12930] = 8'h01;
ROM_MEM[12931] = 8'h04;
ROM_MEM[12932] = 8'h01;
ROM_MEM[12933] = 8'hA5;
ROM_MEM[12934] = 8'hFF;
ROM_MEM[12935] = 8'h01;
ROM_MEM[12936] = 8'h15;
ROM_MEM[12937] = 8'hA1;
ROM_MEM[12938] = 8'h00;
ROM_MEM[12939] = 8'h00;
ROM_MEM[12940] = 8'h02;
ROM_MEM[12941] = 8'h92;
ROM_MEM[12942] = 8'h09;
ROM_MEM[12943] = 8'h00;
ROM_MEM[12944] = 8'h01;
ROM_MEM[12945] = 8'h1E;
ROM_MEM[12946] = 8'h09;
ROM_MEM[12947] = 8'h00;
ROM_MEM[12948] = 8'h01;
ROM_MEM[12949] = 8'h0D;
ROM_MEM[12950] = 8'h09;
ROM_MEM[12951] = 8'h00;
ROM_MEM[12952] = 8'h01;
ROM_MEM[12953] = 8'h03;
ROM_MEM[12954] = 8'h18;
ROM_MEM[12955] = 8'h00;
ROM_MEM[12956] = 8'h02;
ROM_MEM[12957] = 8'h06;
ROM_MEM[12958] = 8'h1C;
ROM_MEM[12959] = 8'hFC;
ROM_MEM[12960] = 8'h01;
ROM_MEM[12961] = 8'h0D;
ROM_MEM[12962] = 8'h06;
ROM_MEM[12963] = 8'h00;
ROM_MEM[12964] = 8'h01;
ROM_MEM[12965] = 8'h18;
ROM_MEM[12966] = 8'h09;
ROM_MEM[12967] = 8'h00;
ROM_MEM[12968] = 8'h01;
ROM_MEM[12969] = 8'h0C;
ROM_MEM[12970] = 8'h0A;
ROM_MEM[12971] = 8'h00;
ROM_MEM[12972] = 8'h02;
ROM_MEM[12973] = 8'h92;
ROM_MEM[12974] = 8'hA0;
ROM_MEM[12975] = 8'h00;
ROM_MEM[12976] = 8'h01;
ROM_MEM[12977] = 8'h1E;
ROM_MEM[12978] = 8'hA0;
ROM_MEM[12979] = 8'h00;
ROM_MEM[12980] = 8'h01;
ROM_MEM[12981] = 8'h09;
ROM_MEM[12982] = 8'hAA;
ROM_MEM[12983] = 8'h00;
ROM_MEM[12984] = 8'h01;
ROM_MEM[12985] = 8'h04;
ROM_MEM[12986] = 8'hA0;
ROM_MEM[12987] = 8'h00;
ROM_MEM[12988] = 8'h01;
ROM_MEM[12989] = 8'h13;
ROM_MEM[12990] = 8'hAA;
ROM_MEM[12991] = 8'h00;
ROM_MEM[12992] = 8'h01;
ROM_MEM[12993] = 8'h09;
ROM_MEM[12994] = 8'hA0;
ROM_MEM[12995] = 8'h00;
ROM_MEM[12996] = 8'h01;
ROM_MEM[12997] = 8'h0A;
ROM_MEM[12998] = 8'hAA;
ROM_MEM[12999] = 8'h00;
ROM_MEM[13000] = 8'h01;
ROM_MEM[13001] = 8'h0E;
ROM_MEM[13002] = 8'hA0;
ROM_MEM[13003] = 8'h00;
ROM_MEM[13004] = 8'h01;
ROM_MEM[13005] = 8'h0C;
ROM_MEM[13006] = 8'hAA;
ROM_MEM[13007] = 8'h00;
ROM_MEM[13008] = 8'h00;
ROM_MEM[13009] = 8'h08;
ROM_MEM[13010] = 8'h6D;
ROM_MEM[13011] = 8'h08;
ROM_MEM[13012] = 8'h6D;
ROM_MEM[13013] = 8'h70;
ROM_MEM[13014] = 8'h08;
ROM_MEM[13015] = 8'h6E;
ROM_MEM[13016] = 8'h0D;
ROM_MEM[13017] = 8'h6E;
ROM_MEM[13018] = 8'hAD;
ROM_MEM[13019] = 8'h06;
ROM_MEM[13020] = 8'h68;
ROM_MEM[13021] = 8'h59;
ROM_MEM[13022] = 8'h68;
ROM_MEM[13023] = 8'h79;
ROM_MEM[13024] = 8'h68;
ROM_MEM[13025] = 8'hAE;
ROM_MEM[13026] = 8'h68;
ROM_MEM[13027] = 8'hD6;
ROM_MEM[13028] = 8'h06;
ROM_MEM[13029] = 8'h68;
ROM_MEM[13030] = 8'hAD;
ROM_MEM[13031] = 8'h68;
ROM_MEM[13032] = 8'hAD;
ROM_MEM[13033] = 8'h69;
ROM_MEM[13034] = 8'h02;
ROM_MEM[13035] = 8'h69;
ROM_MEM[13036] = 8'h02;
ROM_MEM[13037] = 8'h30;
ROM_MEM[13038] = 8'h69;
ROM_MEM[13039] = 8'h03;
ROM_MEM[13040] = 8'h69;
ROM_MEM[13041] = 8'h1F;
ROM_MEM[13042] = 8'h69;
ROM_MEM[13043] = 8'h7D;
ROM_MEM[13044] = 8'h69;
ROM_MEM[13045] = 8'h8D;
ROM_MEM[13046] = 8'h05;
ROM_MEM[13047] = 8'h69;
ROM_MEM[13048] = 8'hF3;
ROM_MEM[13049] = 8'h69;
ROM_MEM[13050] = 8'hF7;
ROM_MEM[13051] = 8'h69;
ROM_MEM[13052] = 8'hF3;
ROM_MEM[13053] = 8'h69;
ROM_MEM[13054] = 8'hF7;
ROM_MEM[13055] = 8'h10;
ROM_MEM[13056] = 8'h6A;
ROM_MEM[13057] = 8'h14;
ROM_MEM[13058] = 8'h6A;
ROM_MEM[13059] = 8'h18;
ROM_MEM[13060] = 8'h20;
ROM_MEM[13061] = 8'h6A;
ROM_MEM[13062] = 8'h25;
ROM_MEM[13063] = 8'h6A;
ROM_MEM[13064] = 8'h31;
ROM_MEM[13065] = 8'h08;
ROM_MEM[13066] = 8'h6A;
ROM_MEM[13067] = 8'h5A;
ROM_MEM[13068] = 8'h6A;
ROM_MEM[13069] = 8'h8E;
ROM_MEM[13070] = 8'hFF;
ROM_MEM[13071] = 8'h6A;
ROM_MEM[13072] = 8'hAB;
ROM_MEM[13073] = 8'h6A;
ROM_MEM[13074] = 8'hCB;
ROM_MEM[13075] = 8'h6A;
ROM_MEM[13076] = 8'hAF;
ROM_MEM[13077] = 8'h6A;
ROM_MEM[13078] = 8'hCB;
ROM_MEM[13079] = 8'h6A;
ROM_MEM[13080] = 8'hB3;
ROM_MEM[13081] = 8'h6A;
ROM_MEM[13082] = 8'hCB;
ROM_MEM[13083] = 8'h6A;
ROM_MEM[13084] = 8'hB7;
ROM_MEM[13085] = 8'h6A;
ROM_MEM[13086] = 8'hCB;
ROM_MEM[13087] = 8'h6A;
ROM_MEM[13088] = 8'hBB;
ROM_MEM[13089] = 8'h6A;
ROM_MEM[13090] = 8'hCB;
ROM_MEM[13091] = 8'h6A;
ROM_MEM[13092] = 8'hBF;
ROM_MEM[13093] = 8'h6A;
ROM_MEM[13094] = 8'hCB;
ROM_MEM[13095] = 8'h6A;
ROM_MEM[13096] = 8'hC3;
ROM_MEM[13097] = 8'h6A;
ROM_MEM[13098] = 8'hCB;
ROM_MEM[13099] = 8'h6A;
ROM_MEM[13100] = 8'hC7;
ROM_MEM[13101] = 8'h6A;
ROM_MEM[13102] = 8'hCB;
ROM_MEM[13103] = 8'h25;
ROM_MEM[13104] = 8'h6B;
ROM_MEM[13105] = 8'h10;
ROM_MEM[13106] = 8'h6B;
ROM_MEM[13107] = 8'h18;
ROM_MEM[13108] = 8'h6B;
ROM_MEM[13109] = 8'h14;
ROM_MEM[13110] = 8'h6B;
ROM_MEM[13111] = 8'h18;
ROM_MEM[13112] = 8'h6B;
ROM_MEM[13113] = 8'h10;
ROM_MEM[13114] = 8'h6B;
ROM_MEM[13115] = 8'h18;
ROM_MEM[13116] = 8'h08;
ROM_MEM[13117] = 8'h6F;
ROM_MEM[13118] = 8'h3A;
ROM_MEM[13119] = 8'h70;
ROM_MEM[13120] = 8'h1E;
ROM_MEM[13121] = 8'h08;
ROM_MEM[13122] = 8'h70;
ROM_MEM[13123] = 8'hDF;
ROM_MEM[13124] = 8'h72;
ROM_MEM[13125] = 8'h1F;
ROM_MEM[13126] = 8'h30;
ROM_MEM[13127] = 8'h69;
ROM_MEM[13128] = 8'h17;
ROM_MEM[13129] = 8'h69;
ROM_MEM[13130] = 8'h58;
ROM_MEM[13131] = 8'h69;
ROM_MEM[13132] = 8'h85;
ROM_MEM[13133] = 8'h69;
ROM_MEM[13134] = 8'hC2;
ROM_MEM[13135] = 8'h01;
ROM_MEM[13136] = 8'h6B;
ROM_MEM[13137] = 8'h31;
ROM_MEM[13138] = 8'h6B;
ROM_MEM[13139] = 8'h35;
ROM_MEM[13140] = 8'hC0;
ROM_MEM[13141] = 8'h6B;
ROM_MEM[13142] = 8'h46;
ROM_MEM[13143] = 8'h6B;
ROM_MEM[13144] = 8'h4E;
ROM_MEM[13145] = 8'h6B;
ROM_MEM[13146] = 8'h6B;
ROM_MEM[13147] = 8'h6B;
ROM_MEM[13148] = 8'h73;
ROM_MEM[13149] = 8'hE2;
ROM_MEM[13150] = 8'h6B;
ROM_MEM[13151] = 8'h8C;
ROM_MEM[13152] = 8'h6C;
ROM_MEM[13153] = 8'h00;
ROM_MEM[13154] = 8'h6B;
ROM_MEM[13155] = 8'hAC;
ROM_MEM[13156] = 8'h6C;
ROM_MEM[13157] = 8'h00;
ROM_MEM[13158] = 8'h6B;
ROM_MEM[13159] = 8'hC8;
ROM_MEM[13160] = 8'h6C;
ROM_MEM[13161] = 8'h00;
ROM_MEM[13162] = 8'h6B;
ROM_MEM[13163] = 8'hE4;
ROM_MEM[13164] = 8'h6C;
ROM_MEM[13165] = 8'h00;
ROM_MEM[13166] = 8'h08;
ROM_MEM[13167] = 8'h72;
ROM_MEM[13168] = 8'h8C;
ROM_MEM[13169] = 8'h72;
ROM_MEM[13170] = 8'hAC;
ROM_MEM[13171] = 8'h30;
ROM_MEM[13172] = 8'h6C;
ROM_MEM[13173] = 8'h0D;
ROM_MEM[13174] = 8'h6C;
ROM_MEM[13175] = 8'h2D;
ROM_MEM[13176] = 8'h6C;
ROM_MEM[13177] = 8'h6A;
ROM_MEM[13178] = 8'h6C;
ROM_MEM[13179] = 8'h7A;
ROM_MEM[13180] = 8'h30;
ROM_MEM[13181] = 8'h69;
ROM_MEM[13182] = 8'h57;
ROM_MEM[13183] = 8'h69;
ROM_MEM[13184] = 8'h57;
ROM_MEM[13185] = 8'h69;
ROM_MEM[13186] = 8'hC1;
ROM_MEM[13187] = 8'h69;
ROM_MEM[13188] = 8'hC1;
ROM_MEM[13189] = 8'h80;
ROM_MEM[13190] = 8'h6C;
ROM_MEM[13191] = 8'h9B;
ROM_MEM[13192] = 8'h6C;
ROM_MEM[13193] = 8'hA3;
ROM_MEM[13194] = 8'h80;
ROM_MEM[13195] = 8'h6C;
ROM_MEM[13196] = 8'h9F;
ROM_MEM[13197] = 8'h6C;
ROM_MEM[13198] = 8'hA3;
ROM_MEM[13199] = 8'hFF;
ROM_MEM[13200] = 8'h6C;
ROM_MEM[13201] = 8'hA8;
ROM_MEM[13202] = 8'h6C;
ROM_MEM[13203] = 8'hAC;
ROM_MEM[13204] = 8'h6C;
ROM_MEM[13205] = 8'hB1;
ROM_MEM[13206] = 8'h6C;
ROM_MEM[13207] = 8'hB5;
ROM_MEM[13208] = 8'h6C;
ROM_MEM[13209] = 8'hBA;
ROM_MEM[13210] = 8'h6C;
ROM_MEM[13211] = 8'hBE;
ROM_MEM[13212] = 8'h6C;
ROM_MEM[13213] = 8'hC7;
ROM_MEM[13214] = 8'h6C;
ROM_MEM[13215] = 8'hCB;
ROM_MEM[13216] = 8'h6C;
ROM_MEM[13217] = 8'hA8;
ROM_MEM[13218] = 8'h6C;
ROM_MEM[13219] = 8'hD4;
ROM_MEM[13220] = 8'h6C;
ROM_MEM[13221] = 8'hB1;
ROM_MEM[13222] = 8'h6C;
ROM_MEM[13223] = 8'hE1;
ROM_MEM[13224] = 8'h6C;
ROM_MEM[13225] = 8'hBA;
ROM_MEM[13226] = 8'h6C;
ROM_MEM[13227] = 8'hEE;
ROM_MEM[13228] = 8'h6C;
ROM_MEM[13229] = 8'hC7;
ROM_MEM[13230] = 8'h6C;
ROM_MEM[13231] = 8'hFB;
ROM_MEM[13232] = 8'h10;
ROM_MEM[13233] = 8'h8E;
ROM_MEM[13234] = 8'h72;
ROM_MEM[13235] = 8'hD1;
ROM_MEM[13236] = 8'h7E;
ROM_MEM[13237] = 8'h74;
ROM_MEM[13238] = 8'h43;
ROM_MEM[13239] = 8'h10;
ROM_MEM[13240] = 8'h8E;
ROM_MEM[13241] = 8'h72;
ROM_MEM[13242] = 8'hD6;
ROM_MEM[13243] = 8'h7E;
ROM_MEM[13244] = 8'h74;
ROM_MEM[13245] = 8'h43;
ROM_MEM[13246] = 8'h10;
ROM_MEM[13247] = 8'h8E;
ROM_MEM[13248] = 8'h73;
ROM_MEM[13249] = 8'h54;
ROM_MEM[13250] = 8'h7E;
ROM_MEM[13251] = 8'h74;
ROM_MEM[13252] = 8'h43;
ROM_MEM[13253] = 8'h10;
ROM_MEM[13254] = 8'h8E;
ROM_MEM[13255] = 8'h72;
ROM_MEM[13256] = 8'hED;
ROM_MEM[13257] = 8'h20;
ROM_MEM[13258] = 8'h78;
ROM_MEM[13259] = 8'h10;
ROM_MEM[13260] = 8'h8E;
ROM_MEM[13261] = 8'h73;
ROM_MEM[13262] = 8'h7C;
ROM_MEM[13263] = 8'h20;
ROM_MEM[13264] = 8'h72;
ROM_MEM[13265] = 8'h10;
ROM_MEM[13266] = 8'h8E;
ROM_MEM[13267] = 8'h72;
ROM_MEM[13268] = 8'hF6;
ROM_MEM[13269] = 8'h20;
ROM_MEM[13270] = 8'h6C;
ROM_MEM[13271] = 8'h10;
ROM_MEM[13272] = 8'h8E;
ROM_MEM[13273] = 8'h72;
ROM_MEM[13274] = 8'hFF;
ROM_MEM[13275] = 8'h20;
ROM_MEM[13276] = 8'h66;
ROM_MEM[13277] = 8'h10;
ROM_MEM[13278] = 8'h8E;
ROM_MEM[13279] = 8'h73;
ROM_MEM[13280] = 8'h04;
ROM_MEM[13281] = 8'h20;
ROM_MEM[13282] = 8'h60;
ROM_MEM[13283] = 8'h10;
ROM_MEM[13284] = 8'h8E;
ROM_MEM[13285] = 8'h72;
ROM_MEM[13286] = 8'hDB;
ROM_MEM[13287] = 8'h20;
ROM_MEM[13288] = 8'h5A;
ROM_MEM[13289] = 8'h10;
ROM_MEM[13290] = 8'h8E;
ROM_MEM[13291] = 8'h72;
ROM_MEM[13292] = 8'hE4;
ROM_MEM[13293] = 8'h20;
ROM_MEM[13294] = 8'h54;
ROM_MEM[13295] = 8'h10;
ROM_MEM[13296] = 8'h8E;
ROM_MEM[13297] = 8'h73;
ROM_MEM[13298] = 8'h09;
ROM_MEM[13299] = 8'h20;
ROM_MEM[13300] = 8'h4E;
ROM_MEM[13301] = 8'h10;
ROM_MEM[13302] = 8'h8E;
ROM_MEM[13303] = 8'h73;
ROM_MEM[13304] = 8'h0E;
ROM_MEM[13305] = 8'h20;
ROM_MEM[13306] = 8'h48;
ROM_MEM[13307] = 8'h10;
ROM_MEM[13308] = 8'h8E;
ROM_MEM[13309] = 8'h73;
ROM_MEM[13310] = 8'h46;
ROM_MEM[13311] = 8'h20;
ROM_MEM[13312] = 8'h42;
ROM_MEM[13313] = 8'h10;
ROM_MEM[13314] = 8'h8E;
ROM_MEM[13315] = 8'h73;
ROM_MEM[13316] = 8'h2F;
ROM_MEM[13317] = 8'h20;
ROM_MEM[13318] = 8'h3C;
ROM_MEM[13319] = 8'h10;
ROM_MEM[13320] = 8'h8E;
ROM_MEM[13321] = 8'h73;
ROM_MEM[13322] = 8'h3C;
ROM_MEM[13323] = 8'h20;
ROM_MEM[13324] = 8'h36;
ROM_MEM[13325] = 8'h10;
ROM_MEM[13326] = 8'h8E;
ROM_MEM[13327] = 8'h73;
ROM_MEM[13328] = 8'h41;
ROM_MEM[13329] = 8'h20;
ROM_MEM[13330] = 8'h30;
ROM_MEM[13331] = 8'h10;
ROM_MEM[13332] = 8'h8E;
ROM_MEM[13333] = 8'h73;
ROM_MEM[13334] = 8'h4F;
ROM_MEM[13335] = 8'h20;
ROM_MEM[13336] = 8'h2A;
ROM_MEM[13337] = 8'h10;
ROM_MEM[13338] = 8'h8E;
ROM_MEM[13339] = 8'h73;
ROM_MEM[13340] = 8'h5D;
ROM_MEM[13341] = 8'h7E;
ROM_MEM[13342] = 8'h74;
ROM_MEM[13343] = 8'h43;
ROM_MEM[13344] = 8'h10;
ROM_MEM[13345] = 8'h8E;
ROM_MEM[13346] = 8'h73;
ROM_MEM[13347] = 8'h6E;
ROM_MEM[13348] = 8'h7E;
ROM_MEM[13349] = 8'h74;
ROM_MEM[13350] = 8'h43;
ROM_MEM[13351] = 8'h10;
ROM_MEM[13352] = 8'h8E;
ROM_MEM[13353] = 8'h73;
ROM_MEM[13354] = 8'h73;
ROM_MEM[13355] = 8'h7E;
ROM_MEM[13356] = 8'h74;
ROM_MEM[13357] = 8'h43;
ROM_MEM[13358] = 8'h10;
ROM_MEM[13359] = 8'h8E;
ROM_MEM[13360] = 8'h73;
ROM_MEM[13361] = 8'h85;
ROM_MEM[13362] = 8'h7E;
ROM_MEM[13363] = 8'h74;
ROM_MEM[13364] = 8'h43;
ROM_MEM[13365] = 8'h10;
ROM_MEM[13366] = 8'h8E;
ROM_MEM[13367] = 8'h73;
ROM_MEM[13368] = 8'h8A;
ROM_MEM[13369] = 8'h7E;
ROM_MEM[13370] = 8'h74;
ROM_MEM[13371] = 8'h43;
ROM_MEM[13372] = 8'h10;
ROM_MEM[13373] = 8'h8E;
ROM_MEM[13374] = 8'h73;
ROM_MEM[13375] = 8'h8F;
ROM_MEM[13376] = 8'h7E;
ROM_MEM[13377] = 8'h74;
ROM_MEM[13378] = 8'h43;
ROM_MEM[13379] = 8'hA6;
ROM_MEM[13380] = 8'hA0;
ROM_MEM[13381] = 8'hB7;
ROM_MEM[13382] = 8'h21;
ROM_MEM[13383] = 8'h00;
ROM_MEM[13384] = 8'h8E;
ROM_MEM[13385] = 8'h21;
ROM_MEM[13386] = 8'h01;
ROM_MEM[13387] = 8'h78;
ROM_MEM[13388] = 8'h21;
ROM_MEM[13389] = 8'h00;
ROM_MEM[13390] = 8'h24;
ROM_MEM[13391] = 8'h12;
ROM_MEM[13392] = 8'hEC;
ROM_MEM[13393] = 8'hA1;
ROM_MEM[13394] = 8'hED;
ROM_MEM[13395] = 8'h84;
ROM_MEM[13396] = 8'hEC;
ROM_MEM[13397] = 8'hA1;
ROM_MEM[13398] = 8'hED;
ROM_MEM[13399] = 8'h05;
ROM_MEM[13400] = 8'h86;
ROM_MEM[13401] = 8'h01;
ROM_MEM[13402] = 8'hA7;
ROM_MEM[13403] = 8'h03;
ROM_MEM[13404] = 8'hA7;
ROM_MEM[13405] = 8'h02;
ROM_MEM[13406] = 8'hA7;
ROM_MEM[13407] = 8'h08;
ROM_MEM[13408] = 8'hA7;
ROM_MEM[13409] = 8'h07;
ROM_MEM[13410] = 8'h30;
ROM_MEM[13411] = 8'h0A;
ROM_MEM[13412] = 8'hB6;
ROM_MEM[13413] = 8'h21;
ROM_MEM[13414] = 8'h00;
ROM_MEM[13415] = 8'h26;
ROM_MEM[13416] = 8'hE2;
ROM_MEM[13417] = 8'h39;
ROM_MEM[13418] = 8'h8E;
ROM_MEM[13419] = 8'h21;
ROM_MEM[13420] = 8'h01;
ROM_MEM[13421] = 8'hC6;
ROM_MEM[13422] = 8'h00;
ROM_MEM[13423] = 8'h10;
ROM_MEM[13424] = 8'hAE;
ROM_MEM[13425] = 8'h84;
ROM_MEM[13426] = 8'h27;
ROM_MEM[13427] = 8'h31;
ROM_MEM[13428] = 8'h6A;
ROM_MEM[13429] = 8'h02;
ROM_MEM[13430] = 8'h26;
ROM_MEM[13431] = 8'h2D;
ROM_MEM[13432] = 8'h6A;
ROM_MEM[13433] = 8'h03;
ROM_MEM[13434] = 8'h26;
ROM_MEM[13435] = 8'h17;
ROM_MEM[13436] = 8'h31;
ROM_MEM[13437] = 8'h24;
ROM_MEM[13438] = 8'h10;
ROM_MEM[13439] = 8'hAF;
ROM_MEM[13440] = 8'h84;
ROM_MEM[13441] = 8'hA6;
ROM_MEM[13442] = 8'h3C;
ROM_MEM[13443] = 8'h26;
ROM_MEM[13444] = 8'h06;
ROM_MEM[13445] = 8'hA7;
ROM_MEM[13446] = 8'h84;
ROM_MEM[13447] = 8'hA7;
ROM_MEM[13448] = 8'h01;
ROM_MEM[13449] = 8'h20;
ROM_MEM[13450] = 8'h14;
ROM_MEM[13451] = 8'hA7;
ROM_MEM[13452] = 8'h03;
ROM_MEM[13453] = 8'hA6;
ROM_MEM[13454] = 8'h3E;
ROM_MEM[13455] = 8'hA7;
ROM_MEM[13456] = 8'h04;
ROM_MEM[13457] = 8'h20;
ROM_MEM[13458] = 8'h06;
ROM_MEM[13459] = 8'hA6;
ROM_MEM[13460] = 8'h04;
ROM_MEM[13461] = 8'hAB;
ROM_MEM[13462] = 8'h3F;
ROM_MEM[13463] = 8'hA7;
ROM_MEM[13464] = 8'h04;
ROM_MEM[13465] = 8'hA6;
ROM_MEM[13466] = 8'h3D;
ROM_MEM[13467] = 8'hA7;
ROM_MEM[13468] = 8'h02;
ROM_MEM[13469] = 8'hA6;
ROM_MEM[13470] = 8'h04;
ROM_MEM[13471] = 8'h10;
ROM_MEM[13472] = 8'h8E;
ROM_MEM[13473] = 8'h18;
ROM_MEM[13474] = 8'h00;
ROM_MEM[13475] = 8'hA7;
ROM_MEM[13476] = 8'hA5;
ROM_MEM[13477] = 8'h30;
ROM_MEM[13478] = 8'h05;
ROM_MEM[13479] = 8'h5C;
ROM_MEM[13480] = 8'hC1;
ROM_MEM[13481] = 8'h10;
ROM_MEM[13482] = 8'h25;
ROM_MEM[13483] = 8'hC3;
ROM_MEM[13484] = 8'h39;
ROM_MEM[13485] = 8'h72;
ROM_MEM[13486] = 8'hD1;
ROM_MEM[13487] = 8'h72;
ROM_MEM[13488] = 8'hD6;
ROM_MEM[13489] = 8'h72;
ROM_MEM[13490] = 8'hDB;
ROM_MEM[13491] = 8'h72;
ROM_MEM[13492] = 8'hE4;
ROM_MEM[13493] = 8'h72;
ROM_MEM[13494] = 8'hED;
ROM_MEM[13495] = 8'h72;
ROM_MEM[13496] = 8'hF6;
ROM_MEM[13497] = 8'h72;
ROM_MEM[13498] = 8'hFF;
ROM_MEM[13499] = 8'h73;
ROM_MEM[13500] = 8'h04;
ROM_MEM[13501] = 8'h73;
ROM_MEM[13502] = 8'h09;
ROM_MEM[13503] = 8'h73;
ROM_MEM[13504] = 8'h0E;
ROM_MEM[13505] = 8'h73;
ROM_MEM[13506] = 8'h2F;
ROM_MEM[13507] = 8'h73;
ROM_MEM[13508] = 8'h3C;
ROM_MEM[13509] = 8'h73;
ROM_MEM[13510] = 8'h41;
ROM_MEM[13511] = 8'h73;
ROM_MEM[13512] = 8'h46;
ROM_MEM[13513] = 8'h73;
ROM_MEM[13514] = 8'h4F;
ROM_MEM[13515] = 8'h73;
ROM_MEM[13516] = 8'h54;
ROM_MEM[13517] = 8'h73;
ROM_MEM[13518] = 8'h5D;
ROM_MEM[13519] = 8'h73;
ROM_MEM[13520] = 8'h6E;
ROM_MEM[13521] = 8'h73;
ROM_MEM[13522] = 8'h73;
ROM_MEM[13523] = 8'h73;
ROM_MEM[13524] = 8'h7C;
ROM_MEM[13525] = 8'h73;
ROM_MEM[13526] = 8'h85;
ROM_MEM[13527] = 8'h73;
ROM_MEM[13528] = 8'h8A;
ROM_MEM[13529] = 8'h73;
ROM_MEM[13530] = 8'h8F;
ROM_MEM[13531] = 8'h22;
ROM_MEM[13532] = 8'h00;
ROM_MEM[13533] = 8'h01;
ROM_MEM[13534] = 8'h18;
ROM_MEM[13535] = 8'h18;
ROM_MEM[13536] = 8'h00;
ROM_MEM[13537] = 8'h18;
ROM_MEM[13538] = 8'h18;
ROM_MEM[13539] = 8'h22;
ROM_MEM[13540] = 8'h19;
ROM_MEM[13541] = 8'h02;
ROM_MEM[13542] = 8'h18;
ROM_MEM[13543] = 8'h1C;
ROM_MEM[13544] = 8'h00;
ROM_MEM[13545] = 8'h18;
ROM_MEM[13546] = 8'h1C;
ROM_MEM[13547] = 8'h22;
ROM_MEM[13548] = 8'h32;
ROM_MEM[13549] = 8'h04;
ROM_MEM[13550] = 8'h18;
ROM_MEM[13551] = 8'h10;
ROM_MEM[13552] = 8'h00;
ROM_MEM[13553] = 8'h18;
ROM_MEM[13554] = 8'h10;
ROM_MEM[13555] = 8'h22;
ROM_MEM[13556] = 8'h4B;
ROM_MEM[13557] = 8'h08;
ROM_MEM[13558] = 8'h18;
ROM_MEM[13559] = 8'h14;
ROM_MEM[13560] = 8'h00;
ROM_MEM[13561] = 8'h18;
ROM_MEM[13562] = 8'h14;
ROM_MEM[13563] = 8'h22;
ROM_MEM[13564] = 8'h64;
ROM_MEM[13565] = 8'h10;
ROM_MEM[13566] = 8'h18;
ROM_MEM[13567] = 8'h14;
ROM_MEM[13568] = 8'h08;
ROM_MEM[13569] = 8'h18;
ROM_MEM[13570] = 8'h16;
ROM_MEM[13571] = 8'h22;
ROM_MEM[13572] = 8'h7D;
ROM_MEM[13573] = 8'h20;
ROM_MEM[13574] = 8'h18;
ROM_MEM[13575] = 8'h14;
ROM_MEM[13576] = 8'h18;
ROM_MEM[13577] = 8'h18;
ROM_MEM[13578] = 8'h1A;
ROM_MEM[13579] = 8'h22;
ROM_MEM[13580] = 8'h96;
ROM_MEM[13581] = 8'h40;
ROM_MEM[13582] = 8'h18;
ROM_MEM[13583] = 8'h14;
ROM_MEM[13584] = 8'h38;
ROM_MEM[13585] = 8'h18;
ROM_MEM[13586] = 8'h1E;
ROM_MEM[13587] = 8'h22;
ROM_MEM[13588] = 8'hAF;
ROM_MEM[13589] = 8'h80;
ROM_MEM[13590] = 8'h18;
ROM_MEM[13591] = 8'h14;
ROM_MEM[13592] = 8'h78;
ROM_MEM[13593] = 8'h18;
ROM_MEM[13594] = 8'h12;
ROM_MEM[13595] = 8'hBD;
ROM_MEM[13596] = 8'h77;
ROM_MEM[13597] = 8'h06;
ROM_MEM[13598] = 8'hC6;
ROM_MEM[13599] = 8'h02;
ROM_MEM[13600] = 8'hBD;
ROM_MEM[13601] = 8'h77;
ROM_MEM[13602] = 8'h6B;
ROM_MEM[13603] = 8'hBD;
ROM_MEM[13604] = 8'h77;
ROM_MEM[13605] = 8'h0A;
ROM_MEM[13606] = 8'hC6;
ROM_MEM[13607] = 8'h04;
ROM_MEM[13608] = 8'hBD;
ROM_MEM[13609] = 8'h77;
ROM_MEM[13610] = 8'h6B;
ROM_MEM[13611] = 8'hBD;
ROM_MEM[13612] = 8'h77;
ROM_MEM[13613] = 8'h0E;
ROM_MEM[13614] = 8'hC6;
ROM_MEM[13615] = 8'h06;
ROM_MEM[13616] = 8'hBD;
ROM_MEM[13617] = 8'h77;
ROM_MEM[13618] = 8'h6B;
ROM_MEM[13619] = 8'hBD;
ROM_MEM[13620] = 8'h77;
ROM_MEM[13621] = 8'h12;
ROM_MEM[13622] = 8'hC6;
ROM_MEM[13623] = 8'h08;
ROM_MEM[13624] = 8'hBD;
ROM_MEM[13625] = 8'h77;
ROM_MEM[13626] = 8'h6B;
ROM_MEM[13627] = 8'h39;
ROM_MEM[13628] = 8'hBD;
ROM_MEM[13629] = 8'h77;
ROM_MEM[13630] = 8'h06;
ROM_MEM[13631] = 8'hC6;
ROM_MEM[13632] = 8'h0E;
ROM_MEM[13633] = 8'hBD;
ROM_MEM[13634] = 8'h77;
ROM_MEM[13635] = 8'h6B;
ROM_MEM[13636] = 8'hBD;
ROM_MEM[13637] = 8'h77;
ROM_MEM[13638] = 8'h0A;
ROM_MEM[13639] = 8'hC6;
ROM_MEM[13640] = 8'h10;
ROM_MEM[13641] = 8'hBD;
ROM_MEM[13642] = 8'h77;
ROM_MEM[13643] = 8'h6B;
ROM_MEM[13644] = 8'hBD;
ROM_MEM[13645] = 8'h77;
ROM_MEM[13646] = 8'h0E;
ROM_MEM[13647] = 8'hC6;
ROM_MEM[13648] = 8'h12;
ROM_MEM[13649] = 8'hBD;
ROM_MEM[13650] = 8'h77;
ROM_MEM[13651] = 8'h6B;
ROM_MEM[13652] = 8'hBD;
ROM_MEM[13653] = 8'h77;
ROM_MEM[13654] = 8'h12;
ROM_MEM[13655] = 8'hC6;
ROM_MEM[13656] = 8'h14;
ROM_MEM[13657] = 8'hBD;
ROM_MEM[13658] = 8'h77;
ROM_MEM[13659] = 8'h6B;
ROM_MEM[13660] = 8'h39;
ROM_MEM[13661] = 8'hBD;
ROM_MEM[13662] = 8'h77;
ROM_MEM[13663] = 8'h06;
ROM_MEM[13664] = 8'hC6;
ROM_MEM[13665] = 8'h16;
ROM_MEM[13666] = 8'hBD;
ROM_MEM[13667] = 8'h77;
ROM_MEM[13668] = 8'h6B;
ROM_MEM[13669] = 8'hBD;
ROM_MEM[13670] = 8'h77;
ROM_MEM[13671] = 8'h0A;
ROM_MEM[13672] = 8'hC6;
ROM_MEM[13673] = 8'h18;
ROM_MEM[13674] = 8'hBD;
ROM_MEM[13675] = 8'h77;
ROM_MEM[13676] = 8'h6B;
ROM_MEM[13677] = 8'hBD;
ROM_MEM[13678] = 8'h77;
ROM_MEM[13679] = 8'h0E;
ROM_MEM[13680] = 8'hC6;
ROM_MEM[13681] = 8'h1A;
ROM_MEM[13682] = 8'hBD;
ROM_MEM[13683] = 8'h77;
ROM_MEM[13684] = 8'h6B;
ROM_MEM[13685] = 8'hBD;
ROM_MEM[13686] = 8'h77;
ROM_MEM[13687] = 8'h12;
ROM_MEM[13688] = 8'hC6;
ROM_MEM[13689] = 8'h1C;
ROM_MEM[13690] = 8'hBD;
ROM_MEM[13691] = 8'h77;
ROM_MEM[13692] = 8'h6B;
ROM_MEM[13693] = 8'h39;
ROM_MEM[13694] = 8'hBD;
ROM_MEM[13695] = 8'h77;
ROM_MEM[13696] = 8'h06;
ROM_MEM[13697] = 8'hC6;
ROM_MEM[13698] = 8'h1E;
ROM_MEM[13699] = 8'hBD;
ROM_MEM[13700] = 8'h77;
ROM_MEM[13701] = 8'h6B;
ROM_MEM[13702] = 8'hBD;
ROM_MEM[13703] = 8'h77;
ROM_MEM[13704] = 8'h0A;
ROM_MEM[13705] = 8'hC6;
ROM_MEM[13706] = 8'h20;
ROM_MEM[13707] = 8'hBD;
ROM_MEM[13708] = 8'h77;
ROM_MEM[13709] = 8'h6B;
ROM_MEM[13710] = 8'hBD;
ROM_MEM[13711] = 8'h77;
ROM_MEM[13712] = 8'h0E;
ROM_MEM[13713] = 8'hC6;
ROM_MEM[13714] = 8'h22;
ROM_MEM[13715] = 8'hBD;
ROM_MEM[13716] = 8'h77;
ROM_MEM[13717] = 8'h6B;
ROM_MEM[13718] = 8'hBD;
ROM_MEM[13719] = 8'h77;
ROM_MEM[13720] = 8'h12;
ROM_MEM[13721] = 8'hC6;
ROM_MEM[13722] = 8'h24;
ROM_MEM[13723] = 8'hBD;
ROM_MEM[13724] = 8'h77;
ROM_MEM[13725] = 8'h6B;
ROM_MEM[13726] = 8'h39;
ROM_MEM[13727] = 8'hBD;
ROM_MEM[13728] = 8'h77;
ROM_MEM[13729] = 8'h06;
ROM_MEM[13730] = 8'hC6;
ROM_MEM[13731] = 8'h26;
ROM_MEM[13732] = 8'hBD;
ROM_MEM[13733] = 8'h77;
ROM_MEM[13734] = 8'h6B;
ROM_MEM[13735] = 8'hBD;
ROM_MEM[13736] = 8'h77;
ROM_MEM[13737] = 8'h0A;
ROM_MEM[13738] = 8'hC6;
ROM_MEM[13739] = 8'h28;
ROM_MEM[13740] = 8'hBD;
ROM_MEM[13741] = 8'h77;
ROM_MEM[13742] = 8'h6B;
ROM_MEM[13743] = 8'hBD;
ROM_MEM[13744] = 8'h77;
ROM_MEM[13745] = 8'h0E;
ROM_MEM[13746] = 8'hC6;
ROM_MEM[13747] = 8'h2A;
ROM_MEM[13748] = 8'hBD;
ROM_MEM[13749] = 8'h77;
ROM_MEM[13750] = 8'h6B;
ROM_MEM[13751] = 8'hBD;
ROM_MEM[13752] = 8'h77;
ROM_MEM[13753] = 8'h12;
ROM_MEM[13754] = 8'hC6;
ROM_MEM[13755] = 8'h2C;
ROM_MEM[13756] = 8'hBD;
ROM_MEM[13757] = 8'h77;
ROM_MEM[13758] = 8'h6B;
ROM_MEM[13759] = 8'h39;
ROM_MEM[13760] = 8'hBD;
ROM_MEM[13761] = 8'h77;
ROM_MEM[13762] = 8'h06;
ROM_MEM[13763] = 8'hC6;
ROM_MEM[13764] = 8'h2E;
ROM_MEM[13765] = 8'hBD;
ROM_MEM[13766] = 8'h77;
ROM_MEM[13767] = 8'h6B;
ROM_MEM[13768] = 8'hBD;
ROM_MEM[13769] = 8'h77;
ROM_MEM[13770] = 8'h0A;
ROM_MEM[13771] = 8'hC6;
ROM_MEM[13772] = 8'h30;
ROM_MEM[13773] = 8'hBD;
ROM_MEM[13774] = 8'h77;
ROM_MEM[13775] = 8'h6B;
ROM_MEM[13776] = 8'hBD;
ROM_MEM[13777] = 8'h77;
ROM_MEM[13778] = 8'h0E;
ROM_MEM[13779] = 8'hC6;
ROM_MEM[13780] = 8'h32;
ROM_MEM[13781] = 8'hBD;
ROM_MEM[13782] = 8'h77;
ROM_MEM[13783] = 8'h6B;
ROM_MEM[13784] = 8'hBD;
ROM_MEM[13785] = 8'h77;
ROM_MEM[13786] = 8'h12;
ROM_MEM[13787] = 8'hC6;
ROM_MEM[13788] = 8'h34;
ROM_MEM[13789] = 8'hBD;
ROM_MEM[13790] = 8'h77;
ROM_MEM[13791] = 8'h6B;
ROM_MEM[13792] = 8'h39;
ROM_MEM[13793] = 8'hBD;
ROM_MEM[13794] = 8'h77;
ROM_MEM[13795] = 8'h06;
ROM_MEM[13796] = 8'hC6;
ROM_MEM[13797] = 8'h36;
ROM_MEM[13798] = 8'hBD;
ROM_MEM[13799] = 8'h77;
ROM_MEM[13800] = 8'h6B;
ROM_MEM[13801] = 8'hBD;
ROM_MEM[13802] = 8'h77;
ROM_MEM[13803] = 8'h0A;
ROM_MEM[13804] = 8'hC6;
ROM_MEM[13805] = 8'h38;
ROM_MEM[13806] = 8'hBD;
ROM_MEM[13807] = 8'h77;
ROM_MEM[13808] = 8'h6B;
ROM_MEM[13809] = 8'hBD;
ROM_MEM[13810] = 8'h77;
ROM_MEM[13811] = 8'h0E;
ROM_MEM[13812] = 8'hC6;
ROM_MEM[13813] = 8'h3A;
ROM_MEM[13814] = 8'hBD;
ROM_MEM[13815] = 8'h77;
ROM_MEM[13816] = 8'h6B;
ROM_MEM[13817] = 8'hBD;
ROM_MEM[13818] = 8'h77;
ROM_MEM[13819] = 8'h12;
ROM_MEM[13820] = 8'hC6;
ROM_MEM[13821] = 8'h3C;
ROM_MEM[13822] = 8'hBD;
ROM_MEM[13823] = 8'h77;
ROM_MEM[13824] = 8'h6B;
ROM_MEM[13825] = 8'h39;
ROM_MEM[13826] = 8'hBD;
ROM_MEM[13827] = 8'h77;
ROM_MEM[13828] = 8'h06;
ROM_MEM[13829] = 8'hC6;
ROM_MEM[13830] = 8'h3E;
ROM_MEM[13831] = 8'hBD;
ROM_MEM[13832] = 8'h77;
ROM_MEM[13833] = 8'h6B;
ROM_MEM[13834] = 8'hBD;
ROM_MEM[13835] = 8'h77;
ROM_MEM[13836] = 8'h0A;
ROM_MEM[13837] = 8'hC6;
ROM_MEM[13838] = 8'h40;
ROM_MEM[13839] = 8'hBD;
ROM_MEM[13840] = 8'h77;
ROM_MEM[13841] = 8'h6B;
ROM_MEM[13842] = 8'hBD;
ROM_MEM[13843] = 8'h77;
ROM_MEM[13844] = 8'h0E;
ROM_MEM[13845] = 8'hC6;
ROM_MEM[13846] = 8'h42;
ROM_MEM[13847] = 8'hBD;
ROM_MEM[13848] = 8'h77;
ROM_MEM[13849] = 8'h6B;
ROM_MEM[13850] = 8'hBD;
ROM_MEM[13851] = 8'h77;
ROM_MEM[13852] = 8'h12;
ROM_MEM[13853] = 8'hC6;
ROM_MEM[13854] = 8'h44;
ROM_MEM[13855] = 8'hBD;
ROM_MEM[13856] = 8'h77;
ROM_MEM[13857] = 8'h6B;
ROM_MEM[13858] = 8'h39;
ROM_MEM[13859] = 8'hBD;
ROM_MEM[13860] = 8'h77;
ROM_MEM[13861] = 8'h06;
ROM_MEM[13862] = 8'hC6;
ROM_MEM[13863] = 8'h46;
ROM_MEM[13864] = 8'hBD;
ROM_MEM[13865] = 8'h77;
ROM_MEM[13866] = 8'h6B;
ROM_MEM[13867] = 8'hBD;
ROM_MEM[13868] = 8'h77;
ROM_MEM[13869] = 8'h0A;
ROM_MEM[13870] = 8'hC6;
ROM_MEM[13871] = 8'h48;
ROM_MEM[13872] = 8'hBD;
ROM_MEM[13873] = 8'h77;
ROM_MEM[13874] = 8'h6B;
ROM_MEM[13875] = 8'hBD;
ROM_MEM[13876] = 8'h77;
ROM_MEM[13877] = 8'h0E;
ROM_MEM[13878] = 8'hC6;
ROM_MEM[13879] = 8'h4A;
ROM_MEM[13880] = 8'hBD;
ROM_MEM[13881] = 8'h77;
ROM_MEM[13882] = 8'h6B;
ROM_MEM[13883] = 8'hBD;
ROM_MEM[13884] = 8'h77;
ROM_MEM[13885] = 8'h12;
ROM_MEM[13886] = 8'hC6;
ROM_MEM[13887] = 8'h4C;
ROM_MEM[13888] = 8'hBD;
ROM_MEM[13889] = 8'h77;
ROM_MEM[13890] = 8'h6B;
ROM_MEM[13891] = 8'h39;
ROM_MEM[13892] = 8'hBD;
ROM_MEM[13893] = 8'h77;
ROM_MEM[13894] = 8'h06;
ROM_MEM[13895] = 8'hC6;
ROM_MEM[13896] = 8'h4E;
ROM_MEM[13897] = 8'hBD;
ROM_MEM[13898] = 8'h77;
ROM_MEM[13899] = 8'h6B;
ROM_MEM[13900] = 8'hBD;
ROM_MEM[13901] = 8'h77;
ROM_MEM[13902] = 8'h0A;
ROM_MEM[13903] = 8'hC6;
ROM_MEM[13904] = 8'h50;
ROM_MEM[13905] = 8'hBD;
ROM_MEM[13906] = 8'h77;
ROM_MEM[13907] = 8'h6B;
ROM_MEM[13908] = 8'hBD;
ROM_MEM[13909] = 8'h77;
ROM_MEM[13910] = 8'h0E;
ROM_MEM[13911] = 8'hC6;
ROM_MEM[13912] = 8'h52;
ROM_MEM[13913] = 8'hBD;
ROM_MEM[13914] = 8'h77;
ROM_MEM[13915] = 8'h6B;
ROM_MEM[13916] = 8'hBD;
ROM_MEM[13917] = 8'h77;
ROM_MEM[13918] = 8'h12;
ROM_MEM[13919] = 8'hC6;
ROM_MEM[13920] = 8'h54;
ROM_MEM[13921] = 8'hBD;
ROM_MEM[13922] = 8'h77;
ROM_MEM[13923] = 8'h6B;
ROM_MEM[13924] = 8'h39;
ROM_MEM[13925] = 8'hBD;
ROM_MEM[13926] = 8'h77;
ROM_MEM[13927] = 8'h06;
ROM_MEM[13928] = 8'hC6;
ROM_MEM[13929] = 8'h56;
ROM_MEM[13930] = 8'hBD;
ROM_MEM[13931] = 8'h77;
ROM_MEM[13932] = 8'h6B;
ROM_MEM[13933] = 8'hBD;
ROM_MEM[13934] = 8'h77;
ROM_MEM[13935] = 8'h0A;
ROM_MEM[13936] = 8'hC6;
ROM_MEM[13937] = 8'h58;
ROM_MEM[13938] = 8'hBD;
ROM_MEM[13939] = 8'h77;
ROM_MEM[13940] = 8'h6B;
ROM_MEM[13941] = 8'hBD;
ROM_MEM[13942] = 8'h77;
ROM_MEM[13943] = 8'h0E;
ROM_MEM[13944] = 8'hC6;
ROM_MEM[13945] = 8'h5A;
ROM_MEM[13946] = 8'hBD;
ROM_MEM[13947] = 8'h77;
ROM_MEM[13948] = 8'h6B;
ROM_MEM[13949] = 8'hBD;
ROM_MEM[13950] = 8'h77;
ROM_MEM[13951] = 8'h12;
ROM_MEM[13952] = 8'hC6;
ROM_MEM[13953] = 8'h5C;
ROM_MEM[13954] = 8'hBD;
ROM_MEM[13955] = 8'h77;
ROM_MEM[13956] = 8'h6B;
ROM_MEM[13957] = 8'h39;
ROM_MEM[13958] = 8'hBD;
ROM_MEM[13959] = 8'h77;
ROM_MEM[13960] = 8'h0E;
ROM_MEM[13961] = 8'hC6;
ROM_MEM[13962] = 8'h5E;
ROM_MEM[13963] = 8'hBD;
ROM_MEM[13964] = 8'h77;
ROM_MEM[13965] = 8'h6B;
ROM_MEM[13966] = 8'hBD;
ROM_MEM[13967] = 8'h77;
ROM_MEM[13968] = 8'h12;
ROM_MEM[13969] = 8'hC6;
ROM_MEM[13970] = 8'h60;
ROM_MEM[13971] = 8'hBD;
ROM_MEM[13972] = 8'h77;
ROM_MEM[13973] = 8'h6B;
ROM_MEM[13974] = 8'hBD;
ROM_MEM[13975] = 8'h77;
ROM_MEM[13976] = 8'h06;
ROM_MEM[13977] = 8'hC6;
ROM_MEM[13978] = 8'h62;
ROM_MEM[13979] = 8'hBD;
ROM_MEM[13980] = 8'h77;
ROM_MEM[13981] = 8'h6B;
ROM_MEM[13982] = 8'hBD;
ROM_MEM[13983] = 8'h77;
ROM_MEM[13984] = 8'h0A;
ROM_MEM[13985] = 8'hC6;
ROM_MEM[13986] = 8'h64;
ROM_MEM[13987] = 8'hBD;
ROM_MEM[13988] = 8'h77;
ROM_MEM[13989] = 8'h6B;
ROM_MEM[13990] = 8'h39;
ROM_MEM[13991] = 8'h86;
ROM_MEM[13992] = 8'h00;
ROM_MEM[13993] = 8'hB7;
ROM_MEM[13994] = 8'h18;
ROM_MEM[13995] = 8'h37;
ROM_MEM[13996] = 8'hB7;
ROM_MEM[13997] = 8'h18;
ROM_MEM[13998] = 8'h3F;
ROM_MEM[13999] = 8'h97;
ROM_MEM[14000] = 8'h12;
ROM_MEM[14001] = 8'hBD;
ROM_MEM[14002] = 8'h77;
ROM_MEM[14003] = 8'h06;
ROM_MEM[14004] = 8'hBD;
ROM_MEM[14005] = 8'h77;
ROM_MEM[14006] = 8'h0A;
ROM_MEM[14007] = 8'hBD;
ROM_MEM[14008] = 8'h77;
ROM_MEM[14009] = 8'h0E;
ROM_MEM[14010] = 8'hBD;
ROM_MEM[14011] = 8'h77;
ROM_MEM[14012] = 8'h12;
ROM_MEM[14013] = 8'hBD;
ROM_MEM[14014] = 8'h77;
ROM_MEM[14015] = 8'h16;
ROM_MEM[14016] = 8'hBD;
ROM_MEM[14017] = 8'h77;
ROM_MEM[14018] = 8'h1A;
ROM_MEM[14019] = 8'hBD;
ROM_MEM[14020] = 8'h77;
ROM_MEM[14021] = 8'h1E;
ROM_MEM[14022] = 8'hBD;
ROM_MEM[14023] = 8'h77;
ROM_MEM[14024] = 8'h22;
ROM_MEM[14025] = 8'h86;
ROM_MEM[14026] = 8'h03;
ROM_MEM[14027] = 8'hB7;
ROM_MEM[14028] = 8'h18;
ROM_MEM[14029] = 8'h37;
ROM_MEM[14030] = 8'hB7;
ROM_MEM[14031] = 8'h18;
ROM_MEM[14032] = 8'h3F;
ROM_MEM[14033] = 8'h86;
ROM_MEM[14034] = 8'h78;
ROM_MEM[14035] = 8'hB7;
ROM_MEM[14036] = 8'h18;
ROM_MEM[14037] = 8'h30;
ROM_MEM[14038] = 8'h86;
ROM_MEM[14039] = 8'h78;
ROM_MEM[14040] = 8'hB7;
ROM_MEM[14041] = 8'h18;
ROM_MEM[14042] = 8'h38;
ROM_MEM[14043] = 8'h39;
ROM_MEM[14044] = 8'h86;
ROM_MEM[14045] = 8'h00;
ROM_MEM[14046] = 8'hB7;
ROM_MEM[14047] = 8'h18;
ROM_MEM[14048] = 8'h30;
ROM_MEM[14049] = 8'hB7;
ROM_MEM[14050] = 8'h18;
ROM_MEM[14051] = 8'h38;
ROM_MEM[14052] = 8'h86;
ROM_MEM[14053] = 8'h01;
ROM_MEM[14054] = 8'h26;
ROM_MEM[14055] = 8'h0B;
ROM_MEM[14056] = 8'h86;
ROM_MEM[14057] = 8'h78;
ROM_MEM[14058] = 8'hB7;
ROM_MEM[14059] = 8'h18;
ROM_MEM[14060] = 8'h30;
ROM_MEM[14061] = 8'h86;
ROM_MEM[14062] = 8'h78;
ROM_MEM[14063] = 8'hB7;
ROM_MEM[14064] = 8'h18;
ROM_MEM[14065] = 8'h38;
ROM_MEM[14066] = 8'h4F;
ROM_MEM[14067] = 8'h97;
ROM_MEM[14068] = 8'h12;
ROM_MEM[14069] = 8'h8D;
ROM_MEM[14070] = 8'h0F;
ROM_MEM[14071] = 8'h8D;
ROM_MEM[14072] = 8'h11;
ROM_MEM[14073] = 8'h8D;
ROM_MEM[14074] = 8'h13;
ROM_MEM[14075] = 8'h8D;
ROM_MEM[14076] = 8'h15;
ROM_MEM[14077] = 8'h8D;
ROM_MEM[14078] = 8'h17;
ROM_MEM[14079] = 8'h8D;
ROM_MEM[14080] = 8'h19;
ROM_MEM[14081] = 8'h8D;
ROM_MEM[14082] = 8'h1B;
ROM_MEM[14083] = 8'h8D;
ROM_MEM[14084] = 8'h1D;
ROM_MEM[14085] = 8'h39;
ROM_MEM[14086] = 8'h86;
ROM_MEM[14087] = 8'h00;
ROM_MEM[14088] = 8'h20;
ROM_MEM[14089] = 8'h1C;
ROM_MEM[14090] = 8'h86;
ROM_MEM[14091] = 8'h08;
ROM_MEM[14092] = 8'h20;
ROM_MEM[14093] = 8'h18;
ROM_MEM[14094] = 8'h86;
ROM_MEM[14095] = 8'h10;
ROM_MEM[14096] = 8'h20;
ROM_MEM[14097] = 8'h14;
ROM_MEM[14098] = 8'h86;
ROM_MEM[14099] = 8'h18;
ROM_MEM[14100] = 8'h20;
ROM_MEM[14101] = 8'h10;
ROM_MEM[14102] = 8'h86;
ROM_MEM[14103] = 8'h20;
ROM_MEM[14104] = 8'h20;
ROM_MEM[14105] = 8'h0C;
ROM_MEM[14106] = 8'h86;
ROM_MEM[14107] = 8'h28;
ROM_MEM[14108] = 8'h20;
ROM_MEM[14109] = 8'h08;
ROM_MEM[14110] = 8'h86;
ROM_MEM[14111] = 8'h30;
ROM_MEM[14112] = 8'h20;
ROM_MEM[14113] = 8'h04;
ROM_MEM[14114] = 8'h86;
ROM_MEM[14115] = 8'h38;
ROM_MEM[14116] = 8'h20;
ROM_MEM[14117] = 8'h00;
ROM_MEM[14118] = 8'h8E;
ROM_MEM[14119] = 8'h74;
ROM_MEM[14120] = 8'hDB;
ROM_MEM[14121] = 8'h31;
ROM_MEM[14122] = 8'h86;
ROM_MEM[14123] = 8'hEE;
ROM_MEM[14124] = 8'hA4;
ROM_MEM[14125] = 8'hA6;
ROM_MEM[14126] = 8'h22;
ROM_MEM[14127] = 8'h43;
ROM_MEM[14128] = 8'h94;
ROM_MEM[14129] = 8'h11;
ROM_MEM[14130] = 8'h97;
ROM_MEM[14131] = 8'h11;
ROM_MEM[14132] = 8'h86;
ROM_MEM[14133] = 8'h07;
ROM_MEM[14134] = 8'hA7;
ROM_MEM[14135] = 8'h4A;
ROM_MEM[14136] = 8'h86;
ROM_MEM[14137] = 8'hC0;
ROM_MEM[14138] = 8'hA7;
ROM_MEM[14139] = 8'h4C;
ROM_MEM[14140] = 8'h86;
ROM_MEM[14141] = 8'hA0;
ROM_MEM[14142] = 8'hA7;
ROM_MEM[14143] = 8'h4E;
ROM_MEM[14144] = 8'hCC;
ROM_MEM[14145] = 8'h00;
ROM_MEM[14146] = 8'h00;
ROM_MEM[14147] = 8'hED;
ROM_MEM[14148] = 8'hC4;
ROM_MEM[14149] = 8'hA7;
ROM_MEM[14150] = 8'h4D;
ROM_MEM[14151] = 8'hA7;
ROM_MEM[14152] = 8'h4B;
ROM_MEM[14153] = 8'hED;
ROM_MEM[14154] = 8'h48;
ROM_MEM[14155] = 8'hA7;
ROM_MEM[14156] = 8'hC8;
ROM_MEM[14157] = 8'h16;
ROM_MEM[14158] = 8'hED;
ROM_MEM[14159] = 8'hC8;
ROM_MEM[14160] = 8'h12;
ROM_MEM[14161] = 8'hA7;
ROM_MEM[14162] = 8'h4F;
ROM_MEM[14163] = 8'hED;
ROM_MEM[14164] = 8'hC8;
ROM_MEM[14165] = 8'h10;
ROM_MEM[14166] = 8'hFC;
ROM_MEM[14167] = 8'h7A;
ROM_MEM[14168] = 8'h17;
ROM_MEM[14169] = 8'hED;
ROM_MEM[14170] = 8'h42;
ROM_MEM[14171] = 8'hED;
ROM_MEM[14172] = 8'h44;
ROM_MEM[14173] = 8'hAE;
ROM_MEM[14174] = 8'h23;
ROM_MEM[14175] = 8'hD6;
ROM_MEM[14176] = 8'h12;
ROM_MEM[14177] = 8'h27;
ROM_MEM[14178] = 8'h05;
ROM_MEM[14179] = 8'hAE;
ROM_MEM[14180] = 8'h26;
ROM_MEM[14181] = 8'h6F;
ROM_MEM[14182] = 8'h01;
ROM_MEM[14183] = 8'h39;
ROM_MEM[14184] = 8'h6F;
ROM_MEM[14185] = 8'h03;
ROM_MEM[14186] = 8'h39;
ROM_MEM[14187] = 8'h8E;
ROM_MEM[14188] = 8'h58;
ROM_MEM[14189] = 8'hE5;
ROM_MEM[14190] = 8'h3A;
ROM_MEM[14191] = 8'hEC;
ROM_MEM[14192] = 8'h84;
ROM_MEM[14193] = 8'hAE;
ROM_MEM[14194] = 8'hA4;
ROM_MEM[14195] = 8'hED;
ROM_MEM[14196] = 8'h84;
ROM_MEM[14197] = 8'h96;
ROM_MEM[14198] = 8'h11;
ROM_MEM[14199] = 8'hAA;
ROM_MEM[14200] = 8'h22;
ROM_MEM[14201] = 8'h97;
ROM_MEM[14202] = 8'h11;
ROM_MEM[14203] = 8'h39;
ROM_MEM[14204] = 8'h96;
ROM_MEM[14205] = 8'h0A;
ROM_MEM[14206] = 8'h44;
ROM_MEM[14207] = 8'h24;
ROM_MEM[14208] = 8'h11;
ROM_MEM[14209] = 8'h86;
ROM_MEM[14210] = 8'h00;
ROM_MEM[14211] = 8'h8D;
ROM_MEM[14212] = 8'h1E;
ROM_MEM[14213] = 8'h86;
ROM_MEM[14214] = 8'h10;
ROM_MEM[14215] = 8'h8D;
ROM_MEM[14216] = 8'h1A;
ROM_MEM[14217] = 8'h86;
ROM_MEM[14218] = 8'h20;
ROM_MEM[14219] = 8'h8D;
ROM_MEM[14220] = 8'h16;
ROM_MEM[14221] = 8'h86;
ROM_MEM[14222] = 8'h30;
ROM_MEM[14223] = 8'h8D;
ROM_MEM[14224] = 8'h12;
ROM_MEM[14225] = 8'h39;
ROM_MEM[14226] = 8'h86;
ROM_MEM[14227] = 8'h08;
ROM_MEM[14228] = 8'h8D;
ROM_MEM[14229] = 8'h0D;
ROM_MEM[14230] = 8'h86;
ROM_MEM[14231] = 8'h18;
ROM_MEM[14232] = 8'h8D;
ROM_MEM[14233] = 8'h09;
ROM_MEM[14234] = 8'h86;
ROM_MEM[14235] = 8'h28;
ROM_MEM[14236] = 8'h8D;
ROM_MEM[14237] = 8'h05;
ROM_MEM[14238] = 8'h86;
ROM_MEM[14239] = 8'h38;
ROM_MEM[14240] = 8'h8D;
ROM_MEM[14241] = 8'h01;
ROM_MEM[14242] = 8'h39;
ROM_MEM[14243] = 8'h8E;
ROM_MEM[14244] = 8'h74;
ROM_MEM[14245] = 8'hDB;
ROM_MEM[14246] = 8'h31;
ROM_MEM[14247] = 8'h86;
ROM_MEM[14248] = 8'hEE;
ROM_MEM[14249] = 8'hA4;
ROM_MEM[14250] = 8'hA6;
ROM_MEM[14251] = 8'hC4;
ROM_MEM[14252] = 8'h26;
ROM_MEM[14253] = 8'h01;
ROM_MEM[14254] = 8'h39;
ROM_MEM[14255] = 8'h6C;
ROM_MEM[14256] = 8'h4B;
ROM_MEM[14257] = 8'h26;
ROM_MEM[14258] = 8'h02;
ROM_MEM[14259] = 8'h6A;
ROM_MEM[14260] = 8'h4B;
ROM_MEM[14261] = 8'hE6;
ROM_MEM[14262] = 8'h4C;
ROM_MEM[14263] = 8'h86;
ROM_MEM[14264] = 8'hFF;
ROM_MEM[14265] = 8'hE3;
ROM_MEM[14266] = 8'h48;
ROM_MEM[14267] = 8'hED;
ROM_MEM[14268] = 8'h48;
ROM_MEM[14269] = 8'h10;
ROM_MEM[14270] = 8'h2A;
ROM_MEM[14271] = 8'h00;
ROM_MEM[14272] = 8'h65;
ROM_MEM[14273] = 8'hAE;
ROM_MEM[14274] = 8'hC4;
ROM_MEM[14275] = 8'hE6;
ROM_MEM[14276] = 8'h81;
ROM_MEM[14277] = 8'hAF;
ROM_MEM[14278] = 8'hC4;
ROM_MEM[14279] = 8'h5D;
ROM_MEM[14280] = 8'h10;
ROM_MEM[14281] = 8'h2B;
ROM_MEM[14282] = 8'h00;
ROM_MEM[14283] = 8'hCE;
ROM_MEM[14284] = 8'h27;
ROM_MEM[14285] = 8'h02;
ROM_MEM[14286] = 8'hEB;
ROM_MEM[14287] = 8'h4D;
ROM_MEM[14288] = 8'h96;
ROM_MEM[14289] = 8'h12;
ROM_MEM[14290] = 8'h27;
ROM_MEM[14291] = 8'h03;
ROM_MEM[14292] = 8'h4F;
ROM_MEM[14293] = 8'h20;
ROM_MEM[14294] = 8'h0E;
ROM_MEM[14295] = 8'h58;
ROM_MEM[14296] = 8'h8E;
ROM_MEM[14297] = 8'h79;
ROM_MEM[14298] = 8'h53;
ROM_MEM[14299] = 8'h3A;
ROM_MEM[14300] = 8'hEC;
ROM_MEM[14301] = 8'h46;
ROM_MEM[14302] = 8'hA3;
ROM_MEM[14303] = 8'h84;
ROM_MEM[14304] = 8'hED;
ROM_MEM[14305] = 8'hC8;
ROM_MEM[14306] = 8'h10;
ROM_MEM[14307] = 8'hEC;
ROM_MEM[14308] = 8'h84;
ROM_MEM[14309] = 8'hED;
ROM_MEM[14310] = 8'h46;
ROM_MEM[14311] = 8'hAE;
ROM_MEM[14312] = 8'hC4;
ROM_MEM[14313] = 8'hA6;
ROM_MEM[14314] = 8'h1F;
ROM_MEM[14315] = 8'h26;
ROM_MEM[14316] = 8'h12;
ROM_MEM[14317] = 8'hEC;
ROM_MEM[14318] = 8'hC8;
ROM_MEM[14319] = 8'h12;
ROM_MEM[14320] = 8'h10;
ROM_MEM[14321] = 8'h27;
ROM_MEM[14322] = 8'hFF;
ROM_MEM[14323] = 8'h37;
ROM_MEM[14324] = 8'hED;
ROM_MEM[14325] = 8'hC4;
ROM_MEM[14326] = 8'hCC;
ROM_MEM[14327] = 8'h00;
ROM_MEM[14328] = 8'h00;
ROM_MEM[14329] = 8'hED;
ROM_MEM[14330] = 8'hC8;
ROM_MEM[14331] = 8'h12;
ROM_MEM[14332] = 8'h7E;
ROM_MEM[14333] = 8'h77;
ROM_MEM[14334] = 8'hC1;
ROM_MEM[14335] = 8'h5F;
ROM_MEM[14336] = 8'h44;
ROM_MEM[14337] = 8'h44;
ROM_MEM[14338] = 8'h56;
ROM_MEM[14339] = 8'hE3;
ROM_MEM[14340] = 8'h48;
ROM_MEM[14341] = 8'hED;
ROM_MEM[14342] = 8'h48;
ROM_MEM[14343] = 8'hA6;
ROM_MEM[14344] = 8'h1F;
ROM_MEM[14345] = 8'h84;
ROM_MEM[14346] = 8'h01;
ROM_MEM[14347] = 8'h26;
ROM_MEM[14348] = 8'h11;
ROM_MEM[14349] = 8'hA7;
ROM_MEM[14350] = 8'h4B;
ROM_MEM[14351] = 8'h5F;
ROM_MEM[14352] = 8'hED;
ROM_MEM[14353] = 8'hC8;
ROM_MEM[14354] = 8'h10;
ROM_MEM[14355] = 8'h96;
ROM_MEM[14356] = 8'h11;
ROM_MEM[14357] = 8'hA4;
ROM_MEM[14358] = 8'h25;
ROM_MEM[14359] = 8'h27;
ROM_MEM[14360] = 8'h0D;
ROM_MEM[14361] = 8'h96;
ROM_MEM[14362] = 8'h12;
ROM_MEM[14363] = 8'h26;
ROM_MEM[14364] = 8'h09;
ROM_MEM[14365] = 8'h39;
ROM_MEM[14366] = 8'hA6;
ROM_MEM[14367] = 8'h4F;
ROM_MEM[14368] = 8'h26;
ROM_MEM[14369] = 8'h04;
ROM_MEM[14370] = 8'h5F;
ROM_MEM[14371] = 8'hED;
ROM_MEM[14372] = 8'hC8;
ROM_MEM[14373] = 8'h10;
ROM_MEM[14374] = 8'h96;
ROM_MEM[14375] = 8'h11;
ROM_MEM[14376] = 8'hA4;
ROM_MEM[14377] = 8'h25;
ROM_MEM[14378] = 8'h27;
ROM_MEM[14379] = 8'h05;
ROM_MEM[14380] = 8'h96;
ROM_MEM[14381] = 8'h12;
ROM_MEM[14382] = 8'h26;
ROM_MEM[14383] = 8'h01;
ROM_MEM[14384] = 8'h39;
ROM_MEM[14385] = 8'h96;
ROM_MEM[14386] = 8'h0A;
ROM_MEM[14387] = 8'h84;
ROM_MEM[14388] = 8'h06;
ROM_MEM[14389] = 8'h26;
ROM_MEM[14390] = 8'h06;
ROM_MEM[14391] = 8'h67;
ROM_MEM[14392] = 8'hC8;
ROM_MEM[14393] = 8'h10;
ROM_MEM[14394] = 8'h66;
ROM_MEM[14395] = 8'hC8;
ROM_MEM[14396] = 8'h11;
ROM_MEM[14397] = 8'hE6;
ROM_MEM[14398] = 8'h4B;
ROM_MEM[14399] = 8'h54;
ROM_MEM[14400] = 8'hAE;
ROM_MEM[14401] = 8'h44;
ROM_MEM[14402] = 8'h3A;
ROM_MEM[14403] = 8'hE6;
ROM_MEM[14404] = 8'h84;
ROM_MEM[14405] = 8'h1D;
ROM_MEM[14406] = 8'h0D;
ROM_MEM[14407] = 8'h12;
ROM_MEM[14408] = 8'h26;
ROM_MEM[14409] = 8'h06;
ROM_MEM[14410] = 8'h58;
ROM_MEM[14411] = 8'h49;
ROM_MEM[14412] = 8'h58;
ROM_MEM[14413] = 8'h49;
ROM_MEM[14414] = 8'h58;
ROM_MEM[14415] = 8'h49;
ROM_MEM[14416] = 8'hE3;
ROM_MEM[14417] = 8'h46;
ROM_MEM[14418] = 8'hE3;
ROM_MEM[14419] = 8'hC8;
ROM_MEM[14420] = 8'h10;
ROM_MEM[14421] = 8'hAE;
ROM_MEM[14422] = 8'h23;
ROM_MEM[14423] = 8'h0D;
ROM_MEM[14424] = 8'h12;
ROM_MEM[14425] = 8'h27;
ROM_MEM[14426] = 8'h04;
ROM_MEM[14427] = 8'hAE;
ROM_MEM[14428] = 8'h26;
ROM_MEM[14429] = 8'h20;
ROM_MEM[14430] = 8'h02;
ROM_MEM[14431] = 8'hA7;
ROM_MEM[14432] = 8'h02;
ROM_MEM[14433] = 8'hE7;
ROM_MEM[14434] = 8'h84;
ROM_MEM[14435] = 8'hEC;
ROM_MEM[14436] = 8'h46;
ROM_MEM[14437] = 8'h26;
ROM_MEM[14438] = 8'h06;
ROM_MEM[14439] = 8'h86;
ROM_MEM[14440] = 8'hF0;
ROM_MEM[14441] = 8'h97;
ROM_MEM[14442] = 8'h10;
ROM_MEM[14443] = 8'h20;
ROM_MEM[14444] = 8'h04;
ROM_MEM[14445] = 8'h86;
ROM_MEM[14446] = 8'hFF;
ROM_MEM[14447] = 8'h97;
ROM_MEM[14448] = 8'h10;
ROM_MEM[14449] = 8'hE6;
ROM_MEM[14450] = 8'h4B;
ROM_MEM[14451] = 8'hC1;
ROM_MEM[14452] = 8'h1F;
ROM_MEM[14453] = 8'h25;
ROM_MEM[14454] = 8'h02;
ROM_MEM[14455] = 8'hC6;
ROM_MEM[14456] = 8'h1F;
ROM_MEM[14457] = 8'hAE;
ROM_MEM[14458] = 8'h42;
ROM_MEM[14459] = 8'hA6;
ROM_MEM[14460] = 8'h85;
ROM_MEM[14461] = 8'hAB;
ROM_MEM[14462] = 8'h4A;
ROM_MEM[14463] = 8'h2A;
ROM_MEM[14464] = 8'h01;
ROM_MEM[14465] = 8'h4F;
ROM_MEM[14466] = 8'h81;
ROM_MEM[14467] = 8'h10;
ROM_MEM[14468] = 8'h2D;
ROM_MEM[14469] = 8'h02;
ROM_MEM[14470] = 8'h86;
ROM_MEM[14471] = 8'h0F;
ROM_MEM[14472] = 8'hAA;
ROM_MEM[14473] = 8'h4E;
ROM_MEM[14474] = 8'h94;
ROM_MEM[14475] = 8'h10;
ROM_MEM[14476] = 8'hAE;
ROM_MEM[14477] = 8'h23;
ROM_MEM[14478] = 8'hD6;
ROM_MEM[14479] = 8'h12;
ROM_MEM[14480] = 8'h27;
ROM_MEM[14481] = 8'h05;
ROM_MEM[14482] = 8'hAE;
ROM_MEM[14483] = 8'h26;
ROM_MEM[14484] = 8'hA7;
ROM_MEM[14485] = 8'h01;
ROM_MEM[14486] = 8'h39;
ROM_MEM[14487] = 8'hA7;
ROM_MEM[14488] = 8'h03;
ROM_MEM[14489] = 8'h39;
ROM_MEM[14490] = 8'hAE;
ROM_MEM[14491] = 8'hC4;
ROM_MEM[14492] = 8'hA6;
ROM_MEM[14493] = 8'h1F;
ROM_MEM[14494] = 8'h58;
ROM_MEM[14495] = 8'hC1;
ROM_MEM[14496] = 8'h24;
ROM_MEM[14497] = 8'h10;
ROM_MEM[14498] = 8'h24;
ROM_MEM[14499] = 8'hFF;
ROM_MEM[14500] = 8'h1C;
ROM_MEM[14501] = 8'h8E;
ROM_MEM[14502] = 8'h78;
ROM_MEM[14503] = 8'hAA;
ROM_MEM[14504] = 8'h6E;
ROM_MEM[14505] = 8'h95;
ROM_MEM[14506] = 8'h78;
ROM_MEM[14507] = 8'hEC;
ROM_MEM[14508] = 8'h78;
ROM_MEM[14509] = 8'hEA;
ROM_MEM[14510] = 8'h78;
ROM_MEM[14511] = 8'hF4;
ROM_MEM[14512] = 8'h78;
ROM_MEM[14513] = 8'hF2;
ROM_MEM[14514] = 8'h78;
ROM_MEM[14515] = 8'hFB;
ROM_MEM[14516] = 8'h78;
ROM_MEM[14517] = 8'hF9;
ROM_MEM[14518] = 8'h78;
ROM_MEM[14519] = 8'hDC;
ROM_MEM[14520] = 8'h78;
ROM_MEM[14521] = 8'hCE;
ROM_MEM[14522] = 8'h77;
ROM_MEM[14523] = 8'hC1;
ROM_MEM[14524] = 8'h77;
ROM_MEM[14525] = 8'hC1;
ROM_MEM[14526] = 8'h79;
ROM_MEM[14527] = 8'h00;
ROM_MEM[14528] = 8'h79;
ROM_MEM[14529] = 8'h05;
ROM_MEM[14530] = 8'h79;
ROM_MEM[14531] = 8'h0B;
ROM_MEM[14532] = 8'h79;
ROM_MEM[14533] = 8'h10;
ROM_MEM[14534] = 8'h79;
ROM_MEM[14535] = 8'h23;
ROM_MEM[14536] = 8'h79;
ROM_MEM[14537] = 8'h2E;
ROM_MEM[14538] = 8'h79;
ROM_MEM[14539] = 8'h3D;
ROM_MEM[14540] = 8'h79;
ROM_MEM[14541] = 8'h4B;
ROM_MEM[14542] = 8'h48;
ROM_MEM[14543] = 8'h1F;
ROM_MEM[14544] = 8'h89;
ROM_MEM[14545] = 8'h8E;
ROM_MEM[14546] = 8'h7A;
ROM_MEM[14547] = 8'h1B;
ROM_MEM[14548] = 8'h3A;
ROM_MEM[14549] = 8'hEC;
ROM_MEM[14550] = 8'h84;
ROM_MEM[14551] = 8'hED;
ROM_MEM[14552] = 8'h42;
ROM_MEM[14553] = 8'h7E;
ROM_MEM[14554] = 8'h77;
ROM_MEM[14555] = 8'hC1;
ROM_MEM[14556] = 8'h48;
ROM_MEM[14557] = 8'h1F;
ROM_MEM[14558] = 8'h89;
ROM_MEM[14559] = 8'h8E;
ROM_MEM[14560] = 8'h7A;
ROM_MEM[14561] = 8'h17;
ROM_MEM[14562] = 8'h3A;
ROM_MEM[14563] = 8'hEC;
ROM_MEM[14564] = 8'h84;
ROM_MEM[14565] = 8'hED;
ROM_MEM[14566] = 8'h44;
ROM_MEM[14567] = 8'h7E;
ROM_MEM[14568] = 8'h77;
ROM_MEM[14569] = 8'hC1;
ROM_MEM[14570] = 8'hA0;
ROM_MEM[14571] = 8'h4C;
ROM_MEM[14572] = 8'h40;
ROM_MEM[14573] = 8'hA7;
ROM_MEM[14574] = 8'h4C;
ROM_MEM[14575] = 8'h7E;
ROM_MEM[14576] = 8'h77;
ROM_MEM[14577] = 8'hC1;
ROM_MEM[14578] = 8'hAB;
ROM_MEM[14579] = 8'h4A;
ROM_MEM[14580] = 8'hA7;
ROM_MEM[14581] = 8'h4A;
ROM_MEM[14582] = 8'h7E;
ROM_MEM[14583] = 8'h77;
ROM_MEM[14584] = 8'hC1;
ROM_MEM[14585] = 8'hAB;
ROM_MEM[14586] = 8'h4D;
ROM_MEM[14587] = 8'hA7;
ROM_MEM[14588] = 8'h4D;
ROM_MEM[14589] = 8'h7E;
ROM_MEM[14590] = 8'h77;
ROM_MEM[14591] = 8'hC1;
ROM_MEM[14592] = 8'hA7;
ROM_MEM[14593] = 8'h4E;
ROM_MEM[14594] = 8'h7E;
ROM_MEM[14595] = 8'h77;
ROM_MEM[14596] = 8'hC1;
ROM_MEM[14597] = 8'hB7;
ROM_MEM[14598] = 8'h18;
ROM_MEM[14599] = 8'h30;
ROM_MEM[14600] = 8'h7E;
ROM_MEM[14601] = 8'h77;
ROM_MEM[14602] = 8'hC1;
ROM_MEM[14603] = 8'hA7;
ROM_MEM[14604] = 8'h4F;
ROM_MEM[14605] = 8'h7E;
ROM_MEM[14606] = 8'h77;
ROM_MEM[14607] = 8'hC1;
ROM_MEM[14608] = 8'h48;
ROM_MEM[14609] = 8'h1F;
ROM_MEM[14610] = 8'h89;
ROM_MEM[14611] = 8'h8E;
ROM_MEM[14612] = 8'h58;
ROM_MEM[14613] = 8'hE5;
ROM_MEM[14614] = 8'h3A;
ROM_MEM[14615] = 8'hEC;
ROM_MEM[14616] = 8'hC4;
ROM_MEM[14617] = 8'hED;
ROM_MEM[14618] = 8'hC8;
ROM_MEM[14619] = 8'h12;
ROM_MEM[14620] = 8'hEC;
ROM_MEM[14621] = 8'h84;
ROM_MEM[14622] = 8'hED;
ROM_MEM[14623] = 8'hC4;
ROM_MEM[14624] = 8'h7E;
ROM_MEM[14625] = 8'h77;
ROM_MEM[14626] = 8'hC1;
ROM_MEM[14627] = 8'hA7;
ROM_MEM[14628] = 8'hC8;
ROM_MEM[14629] = 8'h16;
ROM_MEM[14630] = 8'hEC;
ROM_MEM[14631] = 8'hC4;
ROM_MEM[14632] = 8'hED;
ROM_MEM[14633] = 8'hC8;
ROM_MEM[14634] = 8'h14;
ROM_MEM[14635] = 8'h7E;
ROM_MEM[14636] = 8'h77;
ROM_MEM[14637] = 8'hC1;
ROM_MEM[14638] = 8'h6A;
ROM_MEM[14639] = 8'hC8;
ROM_MEM[14640] = 8'h16;
ROM_MEM[14641] = 8'h10;
ROM_MEM[14642] = 8'h27;
ROM_MEM[14643] = 8'hFE;
ROM_MEM[14644] = 8'h8C;
ROM_MEM[14645] = 8'hEC;
ROM_MEM[14646] = 8'hC8;
ROM_MEM[14647] = 8'h14;
ROM_MEM[14648] = 8'hED;
ROM_MEM[14649] = 8'hC4;
ROM_MEM[14650] = 8'h7E;
ROM_MEM[14651] = 8'h77;
ROM_MEM[14652] = 8'hC1;
ROM_MEM[14653] = 8'hAE;
ROM_MEM[14654] = 8'hC4;
ROM_MEM[14655] = 8'h30;
ROM_MEM[14656] = 8'h01;
ROM_MEM[14657] = 8'hAF;
ROM_MEM[14658] = 8'hC8;
ROM_MEM[14659] = 8'h17;
ROM_MEM[14660] = 8'hEC;
ROM_MEM[14661] = 8'h1E;
ROM_MEM[14662] = 8'hED;
ROM_MEM[14663] = 8'hC4;
ROM_MEM[14664] = 8'h7E;
ROM_MEM[14665] = 8'h77;
ROM_MEM[14666] = 8'hC1;
ROM_MEM[14667] = 8'hEC;
ROM_MEM[14668] = 8'hC8;
ROM_MEM[14669] = 8'h17;
ROM_MEM[14670] = 8'hED;
ROM_MEM[14671] = 8'hC4;
ROM_MEM[14672] = 8'h7E;
ROM_MEM[14673] = 8'h77;
ROM_MEM[14674] = 8'hC1;
ROM_MEM[14675] = 8'h00;
ROM_MEM[14676] = 8'h00;
ROM_MEM[14677] = 8'hB4;
ROM_MEM[14678] = 8'h93;
ROM_MEM[14679] = 8'hAA;
ROM_MEM[14680] = 8'h70;
ROM_MEM[14681] = 8'hA0;
ROM_MEM[14682] = 8'hDF;
ROM_MEM[14683] = 8'h97;
ROM_MEM[14684] = 8'hD7;
ROM_MEM[14685] = 8'h8F;
ROM_MEM[14686] = 8'h51;
ROM_MEM[14687] = 8'h87;
ROM_MEM[14688] = 8'h45;
ROM_MEM[14689] = 8'h7F;
ROM_MEM[14690] = 8'hAD;
ROM_MEM[14691] = 8'h78;
ROM_MEM[14692] = 8'h82;
ROM_MEM[14693] = 8'h71;
ROM_MEM[14694] = 8'hBF;
ROM_MEM[14695] = 8'h6B;
ROM_MEM[14696] = 8'h5C;
ROM_MEM[14697] = 8'h65;
ROM_MEM[14698] = 8'h55;
ROM_MEM[14699] = 8'h5F;
ROM_MEM[14700] = 8'hA5;
ROM_MEM[14701] = 8'h5A;
ROM_MEM[14702] = 8'h46;
ROM_MEM[14703] = 8'h55;
ROM_MEM[14704] = 8'h35;
ROM_MEM[14705] = 8'h50;
ROM_MEM[14706] = 8'h6C;
ROM_MEM[14707] = 8'h4B;
ROM_MEM[14708] = 8'hE8;
ROM_MEM[14709] = 8'h47;
ROM_MEM[14710] = 8'hA5;
ROM_MEM[14711] = 8'h43;
ROM_MEM[14712] = 8'h9F;
ROM_MEM[14713] = 8'h3F;
ROM_MEM[14714] = 8'hD3;
ROM_MEM[14715] = 8'h3C;
ROM_MEM[14716] = 8'h3E;
ROM_MEM[14717] = 8'h38;
ROM_MEM[14718] = 8'hDC;
ROM_MEM[14719] = 8'h35;
ROM_MEM[14720] = 8'hAA;
ROM_MEM[14721] = 8'h32;
ROM_MEM[14722] = 8'hA7;
ROM_MEM[14723] = 8'h2F;
ROM_MEM[14724] = 8'hCF;
ROM_MEM[14725] = 8'h2D;
ROM_MEM[14726] = 8'h20;
ROM_MEM[14727] = 8'h2A;
ROM_MEM[14728] = 8'h97;
ROM_MEM[14729] = 8'h28;
ROM_MEM[14730] = 8'h32;
ROM_MEM[14731] = 8'h25;
ROM_MEM[14732] = 8'hF1;
ROM_MEM[14733] = 8'h23;
ROM_MEM[14734] = 8'hCF;
ROM_MEM[14735] = 8'h21;
ROM_MEM[14736] = 8'hCC;
ROM_MEM[14737] = 8'h1F;
ROM_MEM[14738] = 8'hE6;
ROM_MEM[14739] = 8'h1E;
ROM_MEM[14740] = 8'h1B;
ROM_MEM[14741] = 8'h1C;
ROM_MEM[14742] = 8'h6A;
ROM_MEM[14743] = 8'h1A;
ROM_MEM[14744] = 8'hD2;
ROM_MEM[14745] = 8'h19;
ROM_MEM[14746] = 8'h50;
ROM_MEM[14747] = 8'h17;
ROM_MEM[14748] = 8'hE4;
ROM_MEM[14749] = 8'h16;
ROM_MEM[14750] = 8'h8C;
ROM_MEM[14751] = 8'h15;
ROM_MEM[14752] = 8'h48;
ROM_MEM[14753] = 8'h14;
ROM_MEM[14754] = 8'h16;
ROM_MEM[14755] = 8'h12;
ROM_MEM[14756] = 8'hF5;
ROM_MEM[14757] = 8'h11;
ROM_MEM[14758] = 8'hE4;
ROM_MEM[14759] = 8'h10;
ROM_MEM[14760] = 8'hE3;
ROM_MEM[14761] = 8'h0F;
ROM_MEM[14762] = 8'hF0;
ROM_MEM[14763] = 8'h0F;
ROM_MEM[14764] = 8'h0A;
ROM_MEM[14765] = 8'h0E;
ROM_MEM[14766] = 8'h32;
ROM_MEM[14767] = 8'h0D;
ROM_MEM[14768] = 8'h65;
ROM_MEM[14769] = 8'h0C;
ROM_MEM[14770] = 8'hA4;
ROM_MEM[14771] = 8'h0B;
ROM_MEM[14772] = 8'hEE;
ROM_MEM[14773] = 8'h0B;
ROM_MEM[14774] = 8'h43;
ROM_MEM[14775] = 8'h0A;
ROM_MEM[14776] = 8'hA0;
ROM_MEM[14777] = 8'h0A;
ROM_MEM[14778] = 8'h07;
ROM_MEM[14779] = 8'h09;
ROM_MEM[14780] = 8'h77;
ROM_MEM[14781] = 8'h08;
ROM_MEM[14782] = 8'hEE;
ROM_MEM[14783] = 8'h08;
ROM_MEM[14784] = 8'h6E;
ROM_MEM[14785] = 8'h07;
ROM_MEM[14786] = 8'hF4;
ROM_MEM[14787] = 8'h07;
ROM_MEM[14788] = 8'h82;
ROM_MEM[14789] = 8'h07;
ROM_MEM[14790] = 8'h15;
ROM_MEM[14791] = 8'h06;
ROM_MEM[14792] = 8'hAF;
ROM_MEM[14793] = 8'h06;
ROM_MEM[14794] = 8'h4F;
ROM_MEM[14795] = 8'h05;
ROM_MEM[14796] = 8'hF4;
ROM_MEM[14797] = 8'h05;
ROM_MEM[14798] = 8'h9E;
ROM_MEM[14799] = 8'h05;
ROM_MEM[14800] = 8'h4D;
ROM_MEM[14801] = 8'h05;
ROM_MEM[14802] = 8'h00;
ROM_MEM[14803] = 8'h04;
ROM_MEM[14804] = 8'hB8;
ROM_MEM[14805] = 8'h04;
ROM_MEM[14806] = 8'h74;
ROM_MEM[14807] = 8'h04;
ROM_MEM[14808] = 8'h33;
ROM_MEM[14809] = 8'h03;
ROM_MEM[14810] = 8'hF7;
ROM_MEM[14811] = 8'h03;
ROM_MEM[14812] = 8'hBD;
ROM_MEM[14813] = 8'h03;
ROM_MEM[14814] = 8'h87;
ROM_MEM[14815] = 8'h03;
ROM_MEM[14816] = 8'h54;
ROM_MEM[14817] = 8'h03;
ROM_MEM[14818] = 8'h24;
ROM_MEM[14819] = 8'h02;
ROM_MEM[14820] = 8'hF6;
ROM_MEM[14821] = 8'h02;
ROM_MEM[14822] = 8'hCB;
ROM_MEM[14823] = 8'h02;
ROM_MEM[14824] = 8'hA3;
ROM_MEM[14825] = 8'h02;
ROM_MEM[14826] = 8'h7D;
ROM_MEM[14827] = 8'h02;
ROM_MEM[14828] = 8'h58;
ROM_MEM[14829] = 8'h02;
ROM_MEM[14830] = 8'h36;
ROM_MEM[14831] = 8'h02;
ROM_MEM[14832] = 8'h16;
ROM_MEM[14833] = 8'h01;
ROM_MEM[14834] = 8'hF8;
ROM_MEM[14835] = 8'h01;
ROM_MEM[14836] = 8'hDB;
ROM_MEM[14837] = 8'h01;
ROM_MEM[14838] = 8'hC0;
ROM_MEM[14839] = 8'h01;
ROM_MEM[14840] = 8'hA7;
ROM_MEM[14841] = 8'h01;
ROM_MEM[14842] = 8'h8E;
ROM_MEM[14843] = 8'h01;
ROM_MEM[14844] = 8'h78;
ROM_MEM[14845] = 8'h01;
ROM_MEM[14846] = 8'h62;
ROM_MEM[14847] = 8'h01;
ROM_MEM[14848] = 8'h4E;
ROM_MEM[14849] = 8'h01;
ROM_MEM[14850] = 8'h3B;
ROM_MEM[14851] = 8'h01;
ROM_MEM[14852] = 8'h29;
ROM_MEM[14853] = 8'h01;
ROM_MEM[14854] = 8'h18;
ROM_MEM[14855] = 8'h01;
ROM_MEM[14856] = 8'h08;
ROM_MEM[14857] = 8'h00;
ROM_MEM[14858] = 8'hF8;
ROM_MEM[14859] = 8'h00;
ROM_MEM[14860] = 8'hEA;
ROM_MEM[14861] = 8'h00;
ROM_MEM[14862] = 8'hDD;
ROM_MEM[14863] = 8'h00;
ROM_MEM[14864] = 8'hD0;
ROM_MEM[14865] = 8'h00;
ROM_MEM[14866] = 8'hC4;
ROM_MEM[14867] = 8'h00;
ROM_MEM[14868] = 8'hB8;
ROM_MEM[14869] = 8'h00;
ROM_MEM[14870] = 8'hAE;
ROM_MEM[14871] = 8'h7A;
ROM_MEM[14872] = 8'h65;
ROM_MEM[14873] = 8'h7A;
ROM_MEM[14874] = 8'h25;
ROM_MEM[14875] = 8'h7A;
ROM_MEM[14876] = 8'h65;
ROM_MEM[14877] = 8'h7A;
ROM_MEM[14878] = 8'hE5;
ROM_MEM[14879] = 8'h7B;
ROM_MEM[14880] = 8'h05;
ROM_MEM[14881] = 8'h7B;
ROM_MEM[14882] = 8'h25;
ROM_MEM[14883] = 8'h7B;
ROM_MEM[14884] = 8'h45;
ROM_MEM[14885] = 8'hFF;
ROM_MEM[14886] = 8'hFF;
ROM_MEM[14887] = 8'hFF;
ROM_MEM[14888] = 8'hFF;
ROM_MEM[14889] = 8'hFF;
ROM_MEM[14890] = 8'hFF;
ROM_MEM[14891] = 8'hFF;
ROM_MEM[14892] = 8'hFF;
ROM_MEM[14893] = 8'hFF;
ROM_MEM[14894] = 8'hFF;
ROM_MEM[14895] = 8'hFF;
ROM_MEM[14896] = 8'hFF;
ROM_MEM[14897] = 8'hFF;
ROM_MEM[14898] = 8'hFF;
ROM_MEM[14899] = 8'hFF;
ROM_MEM[14900] = 8'hFF;
ROM_MEM[14901] = 8'hFF;
ROM_MEM[14902] = 8'hFF;
ROM_MEM[14903] = 8'hFF;
ROM_MEM[14904] = 8'hFF;
ROM_MEM[14905] = 8'hFF;
ROM_MEM[14906] = 8'hFF;
ROM_MEM[14907] = 8'hFF;
ROM_MEM[14908] = 8'hFF;
ROM_MEM[14909] = 8'hFF;
ROM_MEM[14910] = 8'hFF;
ROM_MEM[14911] = 8'hFF;
ROM_MEM[14912] = 8'hFF;
ROM_MEM[14913] = 8'hFF;
ROM_MEM[14914] = 8'hFF;
ROM_MEM[14915] = 8'hFF;
ROM_MEM[14916] = 8'hFF;
ROM_MEM[14917] = 8'hFF;
ROM_MEM[14918] = 8'hFF;
ROM_MEM[14919] = 8'hFF;
ROM_MEM[14920] = 8'hFF;
ROM_MEM[14921] = 8'hFF;
ROM_MEM[14922] = 8'hFF;
ROM_MEM[14923] = 8'hFF;
ROM_MEM[14924] = 8'hFF;
ROM_MEM[14925] = 8'hFF;
ROM_MEM[14926] = 8'hFF;
ROM_MEM[14927] = 8'hFF;
ROM_MEM[14928] = 8'hFF;
ROM_MEM[14929] = 8'hFF;
ROM_MEM[14930] = 8'hFF;
ROM_MEM[14931] = 8'hFF;
ROM_MEM[14932] = 8'hFF;
ROM_MEM[14933] = 8'hFF;
ROM_MEM[14934] = 8'hFF;
ROM_MEM[14935] = 8'hFF;
ROM_MEM[14936] = 8'hFF;
ROM_MEM[14937] = 8'hFF;
ROM_MEM[14938] = 8'hFF;
ROM_MEM[14939] = 8'hFF;
ROM_MEM[14940] = 8'hFF;
ROM_MEM[14941] = 8'hFF;
ROM_MEM[14942] = 8'hFF;
ROM_MEM[14943] = 8'hFF;
ROM_MEM[14944] = 8'hFF;
ROM_MEM[14945] = 8'hFF;
ROM_MEM[14946] = 8'hFF;
ROM_MEM[14947] = 8'hFF;
ROM_MEM[14948] = 8'hFF;
ROM_MEM[14949] = 8'h00;
ROM_MEM[14950] = 8'h00;
ROM_MEM[14951] = 8'h00;
ROM_MEM[14952] = 8'h00;
ROM_MEM[14953] = 8'h00;
ROM_MEM[14954] = 8'h00;
ROM_MEM[14955] = 8'h00;
ROM_MEM[14956] = 8'h00;
ROM_MEM[14957] = 8'h00;
ROM_MEM[14958] = 8'h00;
ROM_MEM[14959] = 8'h00;
ROM_MEM[14960] = 8'h00;
ROM_MEM[14961] = 8'h00;
ROM_MEM[14962] = 8'h00;
ROM_MEM[14963] = 8'h00;
ROM_MEM[14964] = 8'h00;
ROM_MEM[14965] = 8'h00;
ROM_MEM[14966] = 8'h00;
ROM_MEM[14967] = 8'h00;
ROM_MEM[14968] = 8'h00;
ROM_MEM[14969] = 8'h00;
ROM_MEM[14970] = 8'h00;
ROM_MEM[14971] = 8'h00;
ROM_MEM[14972] = 8'h00;
ROM_MEM[14973] = 8'h00;
ROM_MEM[14974] = 8'h00;
ROM_MEM[14975] = 8'h00;
ROM_MEM[14976] = 8'h00;
ROM_MEM[14977] = 8'h00;
ROM_MEM[14978] = 8'h00;
ROM_MEM[14979] = 8'h00;
ROM_MEM[14980] = 8'h00;
ROM_MEM[14981] = 8'h00;
ROM_MEM[14982] = 8'h00;
ROM_MEM[14983] = 8'h00;
ROM_MEM[14984] = 8'h00;
ROM_MEM[14985] = 8'h00;
ROM_MEM[14986] = 8'h00;
ROM_MEM[14987] = 8'h00;
ROM_MEM[14988] = 8'h00;
ROM_MEM[14989] = 8'h00;
ROM_MEM[14990] = 8'h00;
ROM_MEM[14991] = 8'h00;
ROM_MEM[14992] = 8'h00;
ROM_MEM[14993] = 8'h00;
ROM_MEM[14994] = 8'h00;
ROM_MEM[14995] = 8'h00;
ROM_MEM[14996] = 8'h00;
ROM_MEM[14997] = 8'h00;
ROM_MEM[14998] = 8'h00;
ROM_MEM[14999] = 8'h00;
ROM_MEM[15000] = 8'h00;
ROM_MEM[15001] = 8'h00;
ROM_MEM[15002] = 8'h00;
ROM_MEM[15003] = 8'h00;
ROM_MEM[15004] = 8'h00;
ROM_MEM[15005] = 8'h00;
ROM_MEM[15006] = 8'h00;
ROM_MEM[15007] = 8'h00;
ROM_MEM[15008] = 8'h00;
ROM_MEM[15009] = 8'h00;
ROM_MEM[15010] = 8'h00;
ROM_MEM[15011] = 8'h00;
ROM_MEM[15012] = 8'h00;
ROM_MEM[15013] = 8'h00;
ROM_MEM[15014] = 8'h00;
ROM_MEM[15015] = 8'h00;
ROM_MEM[15016] = 8'h00;
ROM_MEM[15017] = 8'h00;
ROM_MEM[15018] = 8'h00;
ROM_MEM[15019] = 8'h00;
ROM_MEM[15020] = 8'h00;
ROM_MEM[15021] = 8'h00;
ROM_MEM[15022] = 8'h00;
ROM_MEM[15023] = 8'h00;
ROM_MEM[15024] = 8'h00;
ROM_MEM[15025] = 8'h00;
ROM_MEM[15026] = 8'h00;
ROM_MEM[15027] = 8'h00;
ROM_MEM[15028] = 8'h00;
ROM_MEM[15029] = 8'h00;
ROM_MEM[15030] = 8'h00;
ROM_MEM[15031] = 8'h00;
ROM_MEM[15032] = 8'h00;
ROM_MEM[15033] = 8'h00;
ROM_MEM[15034] = 8'h00;
ROM_MEM[15035] = 8'h00;
ROM_MEM[15036] = 8'h00;
ROM_MEM[15037] = 8'h00;
ROM_MEM[15038] = 8'h00;
ROM_MEM[15039] = 8'h00;
ROM_MEM[15040] = 8'h00;
ROM_MEM[15041] = 8'h00;
ROM_MEM[15042] = 8'h00;
ROM_MEM[15043] = 8'h00;
ROM_MEM[15044] = 8'h00;
ROM_MEM[15045] = 8'h00;
ROM_MEM[15046] = 8'h00;
ROM_MEM[15047] = 8'h00;
ROM_MEM[15048] = 8'h00;
ROM_MEM[15049] = 8'h00;
ROM_MEM[15050] = 8'h00;
ROM_MEM[15051] = 8'h00;
ROM_MEM[15052] = 8'h00;
ROM_MEM[15053] = 8'h00;
ROM_MEM[15054] = 8'h00;
ROM_MEM[15055] = 8'h00;
ROM_MEM[15056] = 8'h00;
ROM_MEM[15057] = 8'h00;
ROM_MEM[15058] = 8'h00;
ROM_MEM[15059] = 8'h00;
ROM_MEM[15060] = 8'h00;
ROM_MEM[15061] = 8'h00;
ROM_MEM[15062] = 8'h00;
ROM_MEM[15063] = 8'h00;
ROM_MEM[15064] = 8'h00;
ROM_MEM[15065] = 8'h00;
ROM_MEM[15066] = 8'h00;
ROM_MEM[15067] = 8'h00;
ROM_MEM[15068] = 8'h00;
ROM_MEM[15069] = 8'h00;
ROM_MEM[15070] = 8'h00;
ROM_MEM[15071] = 8'h00;
ROM_MEM[15072] = 8'h00;
ROM_MEM[15073] = 8'h00;
ROM_MEM[15074] = 8'h00;
ROM_MEM[15075] = 8'h00;
ROM_MEM[15076] = 8'h00;
ROM_MEM[15077] = 8'h0A;
ROM_MEM[15078] = 8'h09;
ROM_MEM[15079] = 8'h08;
ROM_MEM[15080] = 8'h07;
ROM_MEM[15081] = 8'h06;
ROM_MEM[15082] = 8'h05;
ROM_MEM[15083] = 8'h04;
ROM_MEM[15084] = 8'h03;
ROM_MEM[15085] = 8'h02;
ROM_MEM[15086] = 8'h02;
ROM_MEM[15087] = 8'h01;
ROM_MEM[15088] = 8'h01;
ROM_MEM[15089] = 8'h01;
ROM_MEM[15090] = 8'h01;
ROM_MEM[15091] = 8'h01;
ROM_MEM[15092] = 8'h01;
ROM_MEM[15093] = 8'h00;
ROM_MEM[15094] = 8'h00;
ROM_MEM[15095] = 8'h00;
ROM_MEM[15096] = 8'h00;
ROM_MEM[15097] = 8'h00;
ROM_MEM[15098] = 8'h00;
ROM_MEM[15099] = 8'h00;
ROM_MEM[15100] = 8'hFF;
ROM_MEM[15101] = 8'hFF;
ROM_MEM[15102] = 8'hFF;
ROM_MEM[15103] = 8'hFF;
ROM_MEM[15104] = 8'hFF;
ROM_MEM[15105] = 8'hFF;
ROM_MEM[15106] = 8'hFF;
ROM_MEM[15107] = 8'hFF;
ROM_MEM[15108] = 8'hFE;
ROM_MEM[15109] = 8'h03;
ROM_MEM[15110] = 8'h07;
ROM_MEM[15111] = 8'h07;
ROM_MEM[15112] = 8'h06;
ROM_MEM[15113] = 8'h05;
ROM_MEM[15114] = 8'h05;
ROM_MEM[15115] = 8'h04;
ROM_MEM[15116] = 8'h04;
ROM_MEM[15117] = 8'h04;
ROM_MEM[15118] = 8'h04;
ROM_MEM[15119] = 8'h03;
ROM_MEM[15120] = 8'h03;
ROM_MEM[15121] = 8'h03;
ROM_MEM[15122] = 8'h03;
ROM_MEM[15123] = 8'h03;
ROM_MEM[15124] = 8'h03;
ROM_MEM[15125] = 8'h02;
ROM_MEM[15126] = 8'h02;
ROM_MEM[15127] = 8'h02;
ROM_MEM[15128] = 8'h02;
ROM_MEM[15129] = 8'h02;
ROM_MEM[15130] = 8'h02;
ROM_MEM[15131] = 8'h01;
ROM_MEM[15132] = 8'h01;
ROM_MEM[15133] = 8'h01;
ROM_MEM[15134] = 8'h01;
ROM_MEM[15135] = 8'h01;
ROM_MEM[15136] = 8'h01;
ROM_MEM[15137] = 8'h00;
ROM_MEM[15138] = 8'h00;
ROM_MEM[15139] = 8'h00;
ROM_MEM[15140] = 8'hFF;
ROM_MEM[15141] = 8'h07;
ROM_MEM[15142] = 8'h06;
ROM_MEM[15143] = 8'h05;
ROM_MEM[15144] = 8'h04;
ROM_MEM[15145] = 8'h04;
ROM_MEM[15146] = 8'h03;
ROM_MEM[15147] = 8'h03;
ROM_MEM[15148] = 8'h02;
ROM_MEM[15149] = 8'h02;
ROM_MEM[15150] = 8'h02;
ROM_MEM[15151] = 8'h01;
ROM_MEM[15152] = 8'h01;
ROM_MEM[15153] = 8'h01;
ROM_MEM[15154] = 8'h01;
ROM_MEM[15155] = 8'h00;
ROM_MEM[15156] = 8'h00;
ROM_MEM[15157] = 8'h00;
ROM_MEM[15158] = 8'h00;
ROM_MEM[15159] = 8'h00;
ROM_MEM[15160] = 8'h00;
ROM_MEM[15161] = 8'h00;
ROM_MEM[15162] = 8'h00;
ROM_MEM[15163] = 8'hFF;
ROM_MEM[15164] = 8'hFF;
ROM_MEM[15165] = 8'hFF;
ROM_MEM[15166] = 8'hFF;
ROM_MEM[15167] = 8'hFF;
ROM_MEM[15168] = 8'hFF;
ROM_MEM[15169] = 8'hFF;
ROM_MEM[15170] = 8'hFF;
ROM_MEM[15171] = 8'hFF;
ROM_MEM[15172] = 8'hFF;
ROM_MEM[15173] = 8'h0A;
ROM_MEM[15174] = 8'h09;
ROM_MEM[15175] = 8'h08;
ROM_MEM[15176] = 8'h07;
ROM_MEM[15177] = 8'h06;
ROM_MEM[15178] = 8'h05;
ROM_MEM[15179] = 8'h04;
ROM_MEM[15180] = 8'h04;
ROM_MEM[15181] = 8'h03;
ROM_MEM[15182] = 8'h03;
ROM_MEM[15183] = 8'h03;
ROM_MEM[15184] = 8'h03;
ROM_MEM[15185] = 8'h03;
ROM_MEM[15186] = 8'h03;
ROM_MEM[15187] = 8'h03;
ROM_MEM[15188] = 8'h03;
ROM_MEM[15189] = 8'h02;
ROM_MEM[15190] = 8'h02;
ROM_MEM[15191] = 8'h02;
ROM_MEM[15192] = 8'h02;
ROM_MEM[15193] = 8'h02;
ROM_MEM[15194] = 8'h02;
ROM_MEM[15195] = 8'h02;
ROM_MEM[15196] = 8'h02;
ROM_MEM[15197] = 8'h02;
ROM_MEM[15198] = 8'h02;
ROM_MEM[15199] = 8'h02;
ROM_MEM[15200] = 8'h02;
ROM_MEM[15201] = 8'h02;
ROM_MEM[15202] = 8'h02;
ROM_MEM[15203] = 8'h02;
ROM_MEM[15204] = 8'h02;
ROM_MEM[15205] = 8'hCC;
ROM_MEM[15206] = 8'h7B;
ROM_MEM[15207] = 8'h6B;
ROM_MEM[15208] = 8'h7E;
ROM_MEM[15209] = 8'h7C;
ROM_MEM[15210] = 8'h1E;
ROM_MEM[15211] = 8'h05;
ROM_MEM[15212] = 8'hFF;
ROM_MEM[15213] = 8'hCC;
ROM_MEM[15214] = 8'h7B;
ROM_MEM[15215] = 8'h73;
ROM_MEM[15216] = 8'h7E;
ROM_MEM[15217] = 8'h7C;
ROM_MEM[15218] = 8'h1E;
ROM_MEM[15219] = 8'hFE;
ROM_MEM[15220] = 8'h07;
ROM_MEM[15221] = 8'hFF;
ROM_MEM[15222] = 8'hCC;
ROM_MEM[15223] = 8'h7B;
ROM_MEM[15224] = 8'h7C;
ROM_MEM[15225] = 8'h7E;
ROM_MEM[15226] = 8'h7C;
ROM_MEM[15227] = 8'h1E;
ROM_MEM[15228] = 8'h06;
ROM_MEM[15229] = 8'hFF;
ROM_MEM[15230] = 8'hCC;
ROM_MEM[15231] = 8'h7B;
ROM_MEM[15232] = 8'h84;
ROM_MEM[15233] = 8'h7E;
ROM_MEM[15234] = 8'h7C;
ROM_MEM[15235] = 8'h1E;
ROM_MEM[15236] = 8'h0A;
ROM_MEM[15237] = 8'h03;
ROM_MEM[15238] = 8'h0A;
ROM_MEM[15239] = 8'hFF;
ROM_MEM[15240] = 8'hCC;
ROM_MEM[15241] = 8'h7B;
ROM_MEM[15242] = 8'h8E;
ROM_MEM[15243] = 8'h7E;
ROM_MEM[15244] = 8'h7C;
ROM_MEM[15245] = 8'h1E;
ROM_MEM[15246] = 8'h01;
ROM_MEM[15247] = 8'hFF;
ROM_MEM[15248] = 8'hCC;
ROM_MEM[15249] = 8'h7B;
ROM_MEM[15250] = 8'h96;
ROM_MEM[15251] = 8'h7E;
ROM_MEM[15252] = 8'h7C;
ROM_MEM[15253] = 8'h1E;
ROM_MEM[15254] = 8'h0A;
ROM_MEM[15255] = 8'h04;
ROM_MEM[15256] = 8'h0A;
ROM_MEM[15257] = 8'hFF;
ROM_MEM[15258] = 8'h8E;
ROM_MEM[15259] = 8'h7B;
ROM_MEM[15260] = 8'hA0;
ROM_MEM[15261] = 8'h7E;
ROM_MEM[15262] = 8'h7C;
ROM_MEM[15263] = 8'h31;
ROM_MEM[15264] = 8'h0B;
ROM_MEM[15265] = 8'h08;
ROM_MEM[15266] = 8'hFF;
ROM_MEM[15267] = 8'hCC;
ROM_MEM[15268] = 8'h7B;
ROM_MEM[15269] = 8'hA9;
ROM_MEM[15270] = 8'h7E;
ROM_MEM[15271] = 8'h7C;
ROM_MEM[15272] = 8'h1E;
ROM_MEM[15273] = 8'h02;
ROM_MEM[15274] = 8'hFF;
ROM_MEM[15275] = 8'hCC;
ROM_MEM[15276] = 8'h7B;
ROM_MEM[15277] = 8'hB1;
ROM_MEM[15278] = 8'h7E;
ROM_MEM[15279] = 8'h7C;
ROM_MEM[15280] = 8'h1E;
ROM_MEM[15281] = 8'h10;
ROM_MEM[15282] = 8'hFF;
ROM_MEM[15283] = 8'hCC;
ROM_MEM[15284] = 8'h7B;
ROM_MEM[15285] = 8'hB8;
ROM_MEM[15286] = 8'h20;
ROM_MEM[15287] = 8'h66;
ROM_MEM[15288] = 8'h0F;
ROM_MEM[15289] = 8'hFF;
ROM_MEM[15290] = 8'hCC;
ROM_MEM[15291] = 8'h7B;
ROM_MEM[15292] = 8'hBF;
ROM_MEM[15293] = 8'h20;
ROM_MEM[15294] = 8'h5F;
ROM_MEM[15295] = 8'h0F;
ROM_MEM[15296] = 8'h10;
ROM_MEM[15297] = 8'hFF;
ROM_MEM[15298] = 8'hCC;
ROM_MEM[15299] = 8'h7B;
ROM_MEM[15300] = 8'hC7;
ROM_MEM[15301] = 8'h20;
ROM_MEM[15302] = 8'h57;
ROM_MEM[15303] = 8'h0A;
ROM_MEM[15304] = 8'h0C;
ROM_MEM[15305] = 8'h0A;
ROM_MEM[15306] = 8'hFF;
ROM_MEM[15307] = 8'hCC;
ROM_MEM[15308] = 8'h7B;
ROM_MEM[15309] = 8'hD0;
ROM_MEM[15310] = 8'h20;
ROM_MEM[15311] = 8'h4E;
ROM_MEM[15312] = 8'h0A;
ROM_MEM[15313] = 8'h0E;
ROM_MEM[15314] = 8'h0A;
ROM_MEM[15315] = 8'hFF;
ROM_MEM[15316] = 8'hCC;
ROM_MEM[15317] = 8'h7B;
ROM_MEM[15318] = 8'hD9;
ROM_MEM[15319] = 8'h20;
ROM_MEM[15320] = 8'h45;
ROM_MEM[15321] = 8'h11;
ROM_MEM[15322] = 8'hFF;
ROM_MEM[15323] = 8'h8E;
ROM_MEM[15324] = 8'h7B;
ROM_MEM[15325] = 8'hE0;
ROM_MEM[15326] = 8'h20;
ROM_MEM[15327] = 8'h51;
ROM_MEM[15328] = 8'hFE;
ROM_MEM[15329] = 8'h13;
ROM_MEM[15330] = 8'hFF;
ROM_MEM[15331] = 8'h8E;
ROM_MEM[15332] = 8'h7B;
ROM_MEM[15333] = 8'hE8;
ROM_MEM[15334] = 8'h20;
ROM_MEM[15335] = 8'h49;
ROM_MEM[15336] = 8'hFE;
ROM_MEM[15337] = 8'hFE;
ROM_MEM[15338] = 8'hFE;
ROM_MEM[15339] = 8'hFE;
ROM_MEM[15340] = 8'hFE;
ROM_MEM[15341] = 8'hFE;
ROM_MEM[15342] = 8'hFE;
ROM_MEM[15343] = 8'h14;
ROM_MEM[15344] = 8'hFF;
ROM_MEM[15345] = 8'h8E;
ROM_MEM[15346] = 8'h7B;
ROM_MEM[15347] = 8'hF6;
ROM_MEM[15348] = 8'h20;
ROM_MEM[15349] = 8'h3B;
ROM_MEM[15350] = 8'h16;
ROM_MEM[15351] = 8'hFF;
ROM_MEM[15352] = 8'hCC;
ROM_MEM[15353] = 8'h7B;
ROM_MEM[15354] = 8'hFD;
ROM_MEM[15355] = 8'h20;
ROM_MEM[15356] = 8'h21;
ROM_MEM[15357] = 8'h17;
ROM_MEM[15358] = 8'hFF;
ROM_MEM[15359] = 8'hCC;
ROM_MEM[15360] = 8'h7C;
ROM_MEM[15361] = 8'h04;
ROM_MEM[15362] = 8'h20;
ROM_MEM[15363] = 8'h1A;
ROM_MEM[15364] = 8'h09;
ROM_MEM[15365] = 8'hFF;
ROM_MEM[15366] = 8'h8E;
ROM_MEM[15367] = 8'h7C;
ROM_MEM[15368] = 8'h0B;
ROM_MEM[15369] = 8'h20;
ROM_MEM[15370] = 8'h26;
ROM_MEM[15371] = 8'h0D;
ROM_MEM[15372] = 8'hFF;
ROM_MEM[15373] = 8'h8E;
ROM_MEM[15374] = 8'h7C;
ROM_MEM[15375] = 8'h12;
ROM_MEM[15376] = 8'h20;
ROM_MEM[15377] = 8'h1F;
ROM_MEM[15378] = 8'h12;
ROM_MEM[15379] = 8'hFF;
ROM_MEM[15380] = 8'hCC;
ROM_MEM[15381] = 8'h7C;
ROM_MEM[15382] = 8'h19;
ROM_MEM[15383] = 8'h20;
ROM_MEM[15384] = 8'h05;
ROM_MEM[15385] = 8'h15;
ROM_MEM[15386] = 8'hFF;
ROM_MEM[15387] = 8'hCC;
ROM_MEM[15388] = 8'h00;
ROM_MEM[15389] = 8'h00;
ROM_MEM[15390] = 8'hDD;
ROM_MEM[15391] = 8'h1B;
ROM_MEM[15392] = 8'hD6;
ROM_MEM[15393] = 8'h1E;
ROM_MEM[15394] = 8'h5C;
ROM_MEM[15395] = 8'hC4;
ROM_MEM[15396] = 8'h0F;
ROM_MEM[15397] = 8'hD7;
ROM_MEM[15398] = 8'h1E;
ROM_MEM[15399] = 8'h58;
ROM_MEM[15400] = 8'h8E;
ROM_MEM[15401] = 8'h23;
ROM_MEM[15402] = 8'h00;
ROM_MEM[15403] = 8'h3A;
ROM_MEM[15404] = 8'hDC;
ROM_MEM[15405] = 8'h1B;
ROM_MEM[15406] = 8'hED;
ROM_MEM[15407] = 8'h84;
ROM_MEM[15408] = 8'h39;
ROM_MEM[15409] = 8'hD6;
ROM_MEM[15410] = 8'h1E;
ROM_MEM[15411] = 8'hD1;
ROM_MEM[15412] = 8'h1D;
ROM_MEM[15413] = 8'h26;
ROM_MEM[15414] = 8'h08;
ROM_MEM[15415] = 8'hD6;
ROM_MEM[15416] = 8'h20;
ROM_MEM[15417] = 8'h26;
ROM_MEM[15418] = 8'h04;
ROM_MEM[15419] = 8'h1F;
ROM_MEM[15420] = 8'h10;
ROM_MEM[15421] = 8'h20;
ROM_MEM[15422] = 8'hDF;
ROM_MEM[15423] = 8'h39;
ROM_MEM[15424] = 8'hD6;
ROM_MEM[15425] = 8'h1E;
ROM_MEM[15426] = 8'hD7;
ROM_MEM[15427] = 8'h1D;
ROM_MEM[15428] = 8'h39;
ROM_MEM[15429] = 8'h86;
ROM_MEM[15430] = 8'h00;
ROM_MEM[15431] = 8'h97;
ROM_MEM[15432] = 8'h1D;
ROM_MEM[15433] = 8'h97;
ROM_MEM[15434] = 8'h1E;
ROM_MEM[15435] = 8'h97;
ROM_MEM[15436] = 8'h16;
ROM_MEM[15437] = 8'h86;
ROM_MEM[15438] = 8'hFF;
ROM_MEM[15439] = 8'h97;
ROM_MEM[15440] = 8'h1F;
ROM_MEM[15441] = 8'h96;
ROM_MEM[15442] = 8'h1D;
ROM_MEM[15443] = 8'h84;
ROM_MEM[15444] = 8'h0F;
ROM_MEM[15445] = 8'h97;
ROM_MEM[15446] = 8'h1D;
ROM_MEM[15447] = 8'h96;
ROM_MEM[15448] = 8'h1E;
ROM_MEM[15449] = 8'h84;
ROM_MEM[15450] = 8'h0F;
ROM_MEM[15451] = 8'h97;
ROM_MEM[15452] = 8'h1E;
ROM_MEM[15453] = 8'h39;
ROM_MEM[15454] = 8'h96;
ROM_MEM[15455] = 8'h1F;
ROM_MEM[15456] = 8'h27;
ROM_MEM[15457] = 8'h3A;
ROM_MEM[15458] = 8'h2A;
ROM_MEM[15459] = 8'h1F;
ROM_MEM[15460] = 8'h48;
ROM_MEM[15461] = 8'h2A;
ROM_MEM[15462] = 8'h0C;
ROM_MEM[15463] = 8'h96;
ROM_MEM[15464] = 8'h80;
ROM_MEM[15465] = 8'h8A;
ROM_MEM[15466] = 8'h23;
ROM_MEM[15467] = 8'h97;
ROM_MEM[15468] = 8'h80;
ROM_MEM[15469] = 8'h86;
ROM_MEM[15470] = 8'hFF;
ROM_MEM[15471] = 8'h97;
ROM_MEM[15472] = 8'h82;
ROM_MEM[15473] = 8'h20;
ROM_MEM[15474] = 8'h06;
ROM_MEM[15475] = 8'h96;
ROM_MEM[15476] = 8'h80;
ROM_MEM[15477] = 8'h84;
ROM_MEM[15478] = 8'hDF;
ROM_MEM[15479] = 8'h97;
ROM_MEM[15480] = 8'h80;
ROM_MEM[15481] = 8'h0A;
ROM_MEM[15482] = 8'h1F;
ROM_MEM[15483] = 8'h2B;
ROM_MEM[15484] = 8'h04;
ROM_MEM[15485] = 8'h86;
ROM_MEM[15486] = 8'h28;
ROM_MEM[15487] = 8'h97;
ROM_MEM[15488] = 8'h1F;
ROM_MEM[15489] = 8'h20;
ROM_MEM[15490] = 8'h18;
ROM_MEM[15491] = 8'h96;
ROM_MEM[15492] = 8'h80;
ROM_MEM[15493] = 8'h8A;
ROM_MEM[15494] = 8'h03;
ROM_MEM[15495] = 8'h97;
ROM_MEM[15496] = 8'h80;
ROM_MEM[15497] = 8'h86;
ROM_MEM[15498] = 8'hFF;
ROM_MEM[15499] = 8'h97;
ROM_MEM[15500] = 8'h82;
ROM_MEM[15501] = 8'h96;
ROM_MEM[15502] = 8'h80;
ROM_MEM[15503] = 8'h84;
ROM_MEM[15504] = 8'hFE;
ROM_MEM[15505] = 8'h97;
ROM_MEM[15506] = 8'h80;
ROM_MEM[15507] = 8'h0A;
ROM_MEM[15508] = 8'h1F;
ROM_MEM[15509] = 8'h26;
ROM_MEM[15510] = 8'h04;
ROM_MEM[15511] = 8'h86;
ROM_MEM[15512] = 8'h00;
ROM_MEM[15513] = 8'h97;
ROM_MEM[15514] = 8'h20;
ROM_MEM[15515] = 8'h39;
ROM_MEM[15516] = 8'h96;
ROM_MEM[15517] = 8'h80;
ROM_MEM[15518] = 8'h84;
ROM_MEM[15519] = 8'h04;
ROM_MEM[15520] = 8'h27;
ROM_MEM[15521] = 8'h0F;
ROM_MEM[15522] = 8'h96;
ROM_MEM[15523] = 8'h0A;
ROM_MEM[15524] = 8'h84;
ROM_MEM[15525] = 8'h03;
ROM_MEM[15526] = 8'h26;
ROM_MEM[15527] = 8'h06;
ROM_MEM[15528] = 8'h0C;
ROM_MEM[15529] = 8'h16;
ROM_MEM[15530] = 8'h10;
ROM_MEM[15531] = 8'h2B;
ROM_MEM[15532] = 8'hFF;
ROM_MEM[15533] = 8'h9F;
ROM_MEM[15534] = 8'h7E;
ROM_MEM[15535] = 8'h7D;
ROM_MEM[15536] = 8'h43;
ROM_MEM[15537] = 8'h86;
ROM_MEM[15538] = 8'h00;
ROM_MEM[15539] = 8'h97;
ROM_MEM[15540] = 8'h16;
ROM_MEM[15541] = 8'h96;
ROM_MEM[15542] = 8'h80;
ROM_MEM[15543] = 8'h8A;
ROM_MEM[15544] = 8'h03;
ROM_MEM[15545] = 8'h97;
ROM_MEM[15546] = 8'h80;
ROM_MEM[15547] = 8'h96;
ROM_MEM[15548] = 8'h20;
ROM_MEM[15549] = 8'h26;
ROM_MEM[15550] = 8'h25;
ROM_MEM[15551] = 8'h96;
ROM_MEM[15552] = 8'h15;
ROM_MEM[15553] = 8'h27;
ROM_MEM[15554] = 8'h05;
ROM_MEM[15555] = 8'h0A;
ROM_MEM[15556] = 8'h15;
ROM_MEM[15557] = 8'h7E;
ROM_MEM[15558] = 8'h7D;
ROM_MEM[15559] = 8'h43;
ROM_MEM[15560] = 8'hD6;
ROM_MEM[15561] = 8'h1D;
ROM_MEM[15562] = 8'hD1;
ROM_MEM[15563] = 8'h1E;
ROM_MEM[15564] = 8'h27;
ROM_MEM[15565] = 8'h75;
ROM_MEM[15566] = 8'h5C;
ROM_MEM[15567] = 8'hC4;
ROM_MEM[15568] = 8'h0F;
ROM_MEM[15569] = 8'hD7;
ROM_MEM[15570] = 8'h1D;
ROM_MEM[15571] = 8'h58;
ROM_MEM[15572] = 8'h8E;
ROM_MEM[15573] = 8'h23;
ROM_MEM[15574] = 8'h00;
ROM_MEM[15575] = 8'hEC;
ROM_MEM[15576] = 8'h85;
ROM_MEM[15577] = 8'hDD;
ROM_MEM[15578] = 8'h19;
ROM_MEM[15579] = 8'h10;
ROM_MEM[15580] = 8'h27;
ROM_MEM[15581] = 8'hFF;
ROM_MEM[15582] = 8'h6E;
ROM_MEM[15583] = 8'h86;
ROM_MEM[15584] = 8'h03;
ROM_MEM[15585] = 8'h97;
ROM_MEM[15586] = 8'h20;
ROM_MEM[15587] = 8'h39;
ROM_MEM[15588] = 8'h81;
ROM_MEM[15589] = 8'h02;
ROM_MEM[15590] = 8'h26;
ROM_MEM[15591] = 8'h1B;
ROM_MEM[15592] = 8'h9E;
ROM_MEM[15593] = 8'h13;
ROM_MEM[15594] = 8'hA6;
ROM_MEM[15595] = 8'h80;
ROM_MEM[15596] = 8'h97;
ROM_MEM[15597] = 8'h82;
ROM_MEM[15598] = 8'h96;
ROM_MEM[15599] = 8'h80;
ROM_MEM[15600] = 8'h84;
ROM_MEM[15601] = 8'hFE;
ROM_MEM[15602] = 8'h97;
ROM_MEM[15603] = 8'h80;
ROM_MEM[15604] = 8'h9F;
ROM_MEM[15605] = 8'h13;
ROM_MEM[15606] = 8'h9C;
ROM_MEM[15607] = 8'h17;
ROM_MEM[15608] = 8'h26;
ROM_MEM[15609] = 8'h49;
ROM_MEM[15610] = 8'h86;
ROM_MEM[15611] = 8'h01;
ROM_MEM[15612] = 8'h97;
ROM_MEM[15613] = 8'h20;
ROM_MEM[15614] = 8'h86;
ROM_MEM[15615] = 8'h80;
ROM_MEM[15616] = 8'h97;
ROM_MEM[15617] = 8'h15;
ROM_MEM[15618] = 8'h39;
ROM_MEM[15619] = 8'h25;
ROM_MEM[15620] = 8'h36;
ROM_MEM[15621] = 8'h9E;
ROM_MEM[15622] = 8'h19;
ROM_MEM[15623] = 8'hE6;
ROM_MEM[15624] = 8'h80;
ROM_MEM[15625] = 8'h9F;
ROM_MEM[15626] = 8'h19;
ROM_MEM[15627] = 8'hC1;
ROM_MEM[15628] = 8'hFE;
ROM_MEM[15629] = 8'h25;
ROM_MEM[15630] = 8'h09;
ROM_MEM[15631] = 8'h27;
ROM_MEM[15632] = 8'hE9;
ROM_MEM[15633] = 8'h0F;
ROM_MEM[15634] = 8'h20;
ROM_MEM[15635] = 8'h86;
ROM_MEM[15636] = 8'hFF;
ROM_MEM[15637] = 8'h97;
ROM_MEM[15638] = 8'h15;
ROM_MEM[15639] = 8'h39;
ROM_MEM[15640] = 8'h8E;
ROM_MEM[15641] = 8'h40;
ROM_MEM[15642] = 8'h02;
ROM_MEM[15643] = 8'h3A;
ROM_MEM[15644] = 8'h3A;
ROM_MEM[15645] = 8'h3A;
ROM_MEM[15646] = 8'h3A;
ROM_MEM[15647] = 8'h8C;
ROM_MEM[15648] = 8'h40;
ROM_MEM[15649] = 8'h62;
ROM_MEM[15650] = 8'h10;
ROM_MEM[15651] = 8'h24;
ROM_MEM[15652] = 8'hFF;
ROM_MEM[15653] = 8'h1F;
ROM_MEM[15654] = 8'hEC;
ROM_MEM[15655] = 8'h84;
ROM_MEM[15656] = 8'hDD;
ROM_MEM[15657] = 8'h13;
ROM_MEM[15658] = 8'hEC;
ROM_MEM[15659] = 8'h02;
ROM_MEM[15660] = 8'hDD;
ROM_MEM[15661] = 8'h17;
ROM_MEM[15662] = 8'h86;
ROM_MEM[15663] = 8'h60;
ROM_MEM[15664] = 8'h97;
ROM_MEM[15665] = 8'h82;
ROM_MEM[15666] = 8'h96;
ROM_MEM[15667] = 8'h80;
ROM_MEM[15668] = 8'h84;
ROM_MEM[15669] = 8'hFE;
ROM_MEM[15670] = 8'h97;
ROM_MEM[15671] = 8'h80;
ROM_MEM[15672] = 8'h0A;
ROM_MEM[15673] = 8'h20;
ROM_MEM[15674] = 8'h39;
ROM_MEM[15675] = 8'h0A;
ROM_MEM[15676] = 8'h15;
ROM_MEM[15677] = 8'h26;
ROM_MEM[15678] = 8'h04;
ROM_MEM[15679] = 8'h86;
ROM_MEM[15680] = 8'h03;
ROM_MEM[15681] = 8'h97;
ROM_MEM[15682] = 8'h20;
ROM_MEM[15683] = 8'h39;
ROM_MEM[15684] = 8'h7E;
ROM_MEM[15685] = 8'h7E;
ROM_MEM[15686] = 8'h27;
ROM_MEM[15687] = 8'h1C;
ROM_MEM[15688] = 8'hEF;
ROM_MEM[15689] = 8'h8E;
ROM_MEM[15690] = 8'h01;
ROM_MEM[15691] = 8'h4D;
ROM_MEM[15692] = 8'h96;
ROM_MEM[15693] = 8'h00;
ROM_MEM[15694] = 8'h81;
ROM_MEM[15695] = 8'h3F;
ROM_MEM[15696] = 8'h26;
ROM_MEM[15697] = 8'hF2;
ROM_MEM[15698] = 8'h1F;
ROM_MEM[15699] = 8'hB8;
ROM_MEM[15700] = 8'h81;
ROM_MEM[15701] = 8'h10;
ROM_MEM[15702] = 8'h26;
ROM_MEM[15703] = 8'hEC;
ROM_MEM[15704] = 8'h30;
ROM_MEM[15705] = 8'h1F;
ROM_MEM[15706] = 8'h27;
ROM_MEM[15707] = 8'hE8;
ROM_MEM[15708] = 8'h04;
ROM_MEM[15709] = 8'h0B;
ROM_MEM[15710] = 8'h24;
ROM_MEM[15711] = 8'hEC;
ROM_MEM[15712] = 8'h86;
ROM_MEM[15713] = 8'h5A;
ROM_MEM[15714] = 8'hB7;
ROM_MEM[15715] = 8'h00;
ROM_MEM[15716] = 8'h00;
ROM_MEM[15717] = 8'h0C;
ROM_MEM[15718] = 8'h0A;
ROM_MEM[15719] = 8'h26;
ROM_MEM[15720] = 8'h2C;
ROM_MEM[15721] = 8'h0C;
ROM_MEM[15722] = 8'h09;
ROM_MEM[15723] = 8'h86;
ROM_MEM[15724] = 8'h03;
ROM_MEM[15725] = 8'hD6;
ROM_MEM[15726] = 8'h0E;
ROM_MEM[15727] = 8'hC1;
ROM_MEM[15728] = 8'h03;
ROM_MEM[15729] = 8'h25;
ROM_MEM[15730] = 8'h02;
ROM_MEM[15731] = 8'h86;
ROM_MEM[15732] = 8'h01;
ROM_MEM[15733] = 8'h94;
ROM_MEM[15734] = 8'h09;
ROM_MEM[15735] = 8'h26;
ROM_MEM[15736] = 8'h1C;
ROM_MEM[15737] = 8'h7F;
ROM_MEM[15738] = 8'h10;
ROM_MEM[15739] = 8'h0F;
ROM_MEM[15740] = 8'h96;
ROM_MEM[15741] = 8'h80;
ROM_MEM[15742] = 8'h84;
ROM_MEM[15743] = 8'h10;
ROM_MEM[15744] = 8'h26;
ROM_MEM[15745] = 8'h13;
ROM_MEM[15746] = 8'h7C;
ROM_MEM[15747] = 8'h10;
ROM_MEM[15748] = 8'h0F;
ROM_MEM[15749] = 8'h5C;
ROM_MEM[15750] = 8'hC1;
ROM_MEM[15751] = 8'h3C;
ROM_MEM[15752] = 8'h25;
ROM_MEM[15753] = 8'h02;
ROM_MEM[15754] = 8'hC6;
ROM_MEM[15755] = 8'h01;
ROM_MEM[15756] = 8'hD7;
ROM_MEM[15757] = 8'h0E;
ROM_MEM[15758] = 8'h8E;
ROM_MEM[15759] = 8'h7F;
ROM_MEM[15760] = 8'h61;
ROM_MEM[15761] = 8'h3A;
ROM_MEM[15762] = 8'h3A;
ROM_MEM[15763] = 8'hAD;
ROM_MEM[15764] = 8'h94;
ROM_MEM[15765] = 8'hBD;
ROM_MEM[15766] = 8'h7C;
ROM_MEM[15767] = 8'h5E;
ROM_MEM[15768] = 8'hBD;
ROM_MEM[15769] = 8'h7D;
ROM_MEM[15770] = 8'hD3;
ROM_MEM[15771] = 8'hD6;
ROM_MEM[15772] = 8'h80;
ROM_MEM[15773] = 8'h96;
ROM_MEM[15774] = 8'h15;
ROM_MEM[15775] = 8'h9A;
ROM_MEM[15776] = 8'h20;
ROM_MEM[15777] = 8'h26;
ROM_MEM[15778] = 8'h1B;
ROM_MEM[15779] = 8'h96;
ROM_MEM[15780] = 8'h11;
ROM_MEM[15781] = 8'h26;
ROM_MEM[15782] = 8'h17;
ROM_MEM[15783] = 8'hB6;
ROM_MEM[15784] = 8'h10;
ROM_MEM[15785] = 8'h0F;
ROM_MEM[15786] = 8'h27;
ROM_MEM[15787] = 8'h06;
ROM_MEM[15788] = 8'h96;
ROM_MEM[15789] = 8'h0E;
ROM_MEM[15790] = 8'h81;
ROM_MEM[15791] = 8'h03;
ROM_MEM[15792] = 8'h23;
ROM_MEM[15793] = 8'h0C;
ROM_MEM[15794] = 8'hBE;
ROM_MEM[15795] = 8'h21;
ROM_MEM[15796] = 8'h2E;
ROM_MEM[15797] = 8'h8C;
ROM_MEM[15798] = 8'h6D;
ROM_MEM[15799] = 8'h08;
ROM_MEM[15800] = 8'h24;
ROM_MEM[15801] = 8'h04;
ROM_MEM[15802] = 8'hC4;
ROM_MEM[15803] = 8'hF7;
ROM_MEM[15804] = 8'h20;
ROM_MEM[15805] = 8'h02;
ROM_MEM[15806] = 8'hCA;
ROM_MEM[15807] = 8'h08;
ROM_MEM[15808] = 8'hD7;
ROM_MEM[15809] = 8'h80;
ROM_MEM[15810] = 8'h96;
ROM_MEM[15811] = 8'h0A;
ROM_MEM[15812] = 8'h44;
ROM_MEM[15813] = 8'h25;
ROM_MEM[15814] = 8'h03;
ROM_MEM[15815] = 8'hBD;
ROM_MEM[15816] = 8'h74;
ROM_MEM[15817] = 8'h6A;
ROM_MEM[15818] = 8'hBD;
ROM_MEM[15819] = 8'h77;
ROM_MEM[15820] = 8'h7C;
ROM_MEM[15821] = 8'hBD;
ROM_MEM[15822] = 8'h7C;
ROM_MEM[15823] = 8'h5E;
ROM_MEM[15824] = 8'h7E;
ROM_MEM[15825] = 8'h7D;
ROM_MEM[15826] = 8'h47;
ROM_MEM[15827] = 8'hD6;
ROM_MEM[15828] = 8'h0D;
ROM_MEM[15829] = 8'hD1;
ROM_MEM[15830] = 8'h0C;
ROM_MEM[15831] = 8'h27;
ROM_MEM[15832] = 8'h19;
ROM_MEM[15833] = 8'h5C;
ROM_MEM[15834] = 8'hC4;
ROM_MEM[15835] = 8'h1F;
ROM_MEM[15836] = 8'hD7;
ROM_MEM[15837] = 8'h0D;
ROM_MEM[15838] = 8'h8E;
ROM_MEM[15839] = 8'h20;
ROM_MEM[15840] = 8'h20;
ROM_MEM[15841] = 8'hE6;
ROM_MEM[15842] = 8'h85;
ROM_MEM[15843] = 8'h10;
ROM_MEM[15844] = 8'h27;
ROM_MEM[15845] = 8'h00;
ROM_MEM[15846] = 8'h40;
ROM_MEM[15847] = 8'hC1;
ROM_MEM[15848] = 8'h3C;
ROM_MEM[15849] = 8'h22;
ROM_MEM[15850] = 8'h07;
ROM_MEM[15851] = 8'h8E;
ROM_MEM[15852] = 8'h7F;
ROM_MEM[15853] = 8'h61;
ROM_MEM[15854] = 8'h3A;
ROM_MEM[15855] = 8'h3A;
ROM_MEM[15856] = 8'hAD;
ROM_MEM[15857] = 8'h94;
ROM_MEM[15858] = 8'h39;
ROM_MEM[15859] = 8'hD6;
ROM_MEM[15860] = 8'h0C;
ROM_MEM[15861] = 8'h8E;
ROM_MEM[15862] = 8'h20;
ROM_MEM[15863] = 8'h20;
ROM_MEM[15864] = 8'h96;
ROM_MEM[15865] = 8'h80;
ROM_MEM[15866] = 8'h2A;
ROM_MEM[15867] = 8'h0A;
ROM_MEM[15868] = 8'hB6;
ROM_MEM[15869] = 8'h08;
ROM_MEM[15870] = 8'h00;
ROM_MEM[15871] = 8'h27;
ROM_MEM[15872] = 8'h26;
ROM_MEM[15873] = 8'h5C;
ROM_MEM[15874] = 8'hC4;
ROM_MEM[15875] = 8'h1F;
ROM_MEM[15876] = 8'hA7;
ROM_MEM[15877] = 8'h85;
ROM_MEM[15878] = 8'h96;
ROM_MEM[15879] = 8'h85;
ROM_MEM[15880] = 8'h2A;
ROM_MEM[15881] = 8'h08;
ROM_MEM[15882] = 8'h86;
ROM_MEM[15883] = 8'h06;
ROM_MEM[15884] = 8'h97;
ROM_MEM[15885] = 8'h9F;
ROM_MEM[15886] = 8'h0C;
ROM_MEM[15887] = 8'h0B;
ROM_MEM[15888] = 8'h29;
ROM_MEM[15889] = 8'h15;
ROM_MEM[15890] = 8'h96;
ROM_MEM[15891] = 8'h80;
ROM_MEM[15892] = 8'h2A;
ROM_MEM[15893] = 8'h0E;
ROM_MEM[15894] = 8'h96;
ROM_MEM[15895] = 8'h85;
ROM_MEM[15896] = 8'hB6;
ROM_MEM[15897] = 8'h08;
ROM_MEM[15898] = 8'h00;
ROM_MEM[15899] = 8'h27;
ROM_MEM[15900] = 8'h0A;
ROM_MEM[15901] = 8'h5C;
ROM_MEM[15902] = 8'hC4;
ROM_MEM[15903] = 8'h1F;
ROM_MEM[15904] = 8'hA7;
ROM_MEM[15905] = 8'h85;
ROM_MEM[15906] = 8'h20;
ROM_MEM[15907] = 8'hEE;
ROM_MEM[15908] = 8'hD7;
ROM_MEM[15909] = 8'h0C;
ROM_MEM[15910] = 8'h3B;
ROM_MEM[15911] = 8'h1A;
ROM_MEM[15912] = 8'h10;
ROM_MEM[15913] = 8'hB6;
ROM_MEM[15914] = 8'h08;
ROM_MEM[15915] = 8'h00;
ROM_MEM[15916] = 8'h10;
ROM_MEM[15917] = 8'hCE;
ROM_MEM[15918] = 8'h10;
ROM_MEM[15919] = 8'h7F;
ROM_MEM[15920] = 8'h86;
ROM_MEM[15921] = 8'h10;
ROM_MEM[15922] = 8'h1F;
ROM_MEM[15923] = 8'h8B;
ROM_MEM[15924] = 8'h86;
ROM_MEM[15925] = 8'hFF;
ROM_MEM[15926] = 8'h97;
ROM_MEM[15927] = 8'h83;
ROM_MEM[15928] = 8'h97;
ROM_MEM[15929] = 8'h82;
ROM_MEM[15930] = 8'h97;
ROM_MEM[15931] = 8'h80;
ROM_MEM[15932] = 8'hC6;
ROM_MEM[15933] = 8'h2B;
ROM_MEM[15934] = 8'hD7;
ROM_MEM[15935] = 8'h81;
ROM_MEM[15936] = 8'h8E;
ROM_MEM[15937] = 8'h18;
ROM_MEM[15938] = 8'h00;
ROM_MEM[15939] = 8'hCC;
ROM_MEM[15940] = 8'h00;
ROM_MEM[15941] = 8'h00;
ROM_MEM[15942] = 8'hED;
ROM_MEM[15943] = 8'h81;
ROM_MEM[15944] = 8'h8C;
ROM_MEM[15945] = 8'h18;
ROM_MEM[15946] = 8'h20;
ROM_MEM[15947] = 8'h25;
ROM_MEM[15948] = 8'hF9;
ROM_MEM[15949] = 8'hB6;
ROM_MEM[15950] = 8'h08;
ROM_MEM[15951] = 8'h00;
ROM_MEM[15952] = 8'hB7;
ROM_MEM[15953] = 8'h00;
ROM_MEM[15954] = 8'h00;
ROM_MEM[15955] = 8'h8E;
ROM_MEM[15956] = 8'h20;
ROM_MEM[15957] = 8'h00;
ROM_MEM[15958] = 8'hCC;
ROM_MEM[15959] = 8'h00;
ROM_MEM[15960] = 8'h00;
ROM_MEM[15961] = 8'hED;
ROM_MEM[15962] = 8'h81;
ROM_MEM[15963] = 8'h8C;
ROM_MEM[15964] = 8'h28;
ROM_MEM[15965] = 8'h00;
ROM_MEM[15966] = 8'h25;
ROM_MEM[15967] = 8'hF9;
ROM_MEM[15968] = 8'h8E;
ROM_MEM[15969] = 8'h10;
ROM_MEM[15970] = 8'h00;
ROM_MEM[15971] = 8'hED;
ROM_MEM[15972] = 8'h81;
ROM_MEM[15973] = 8'h8C;
ROM_MEM[15974] = 8'h10;
ROM_MEM[15975] = 8'h80;
ROM_MEM[15976] = 8'h25;
ROM_MEM[15977] = 8'hF9;
ROM_MEM[15978] = 8'hB7;
ROM_MEM[15979] = 8'h18;
ROM_MEM[15980] = 8'h27;
ROM_MEM[15981] = 8'hB7;
ROM_MEM[15982] = 8'h18;
ROM_MEM[15983] = 8'h2F;
ROM_MEM[15984] = 8'hB7;
ROM_MEM[15985] = 8'h18;
ROM_MEM[15986] = 8'h37;
ROM_MEM[15987] = 8'hB7;
ROM_MEM[15988] = 8'h18;
ROM_MEM[15989] = 8'h3F;
ROM_MEM[15990] = 8'hB7;
ROM_MEM[15991] = 8'h18;
ROM_MEM[15992] = 8'h20;
ROM_MEM[15993] = 8'hB7;
ROM_MEM[15994] = 8'h18;
ROM_MEM[15995] = 8'h28;
ROM_MEM[15996] = 8'hB7;
ROM_MEM[15997] = 8'h18;
ROM_MEM[15998] = 8'h30;
ROM_MEM[15999] = 8'hB7;
ROM_MEM[16000] = 8'h18;
ROM_MEM[16001] = 8'h38;
ROM_MEM[16002] = 8'h86;
ROM_MEM[16003] = 8'h07;
ROM_MEM[16004] = 8'hB7;
ROM_MEM[16005] = 8'h18;
ROM_MEM[16006] = 8'h27;
ROM_MEM[16007] = 8'hB7;
ROM_MEM[16008] = 8'h18;
ROM_MEM[16009] = 8'h2F;
ROM_MEM[16010] = 8'hB7;
ROM_MEM[16011] = 8'h18;
ROM_MEM[16012] = 8'h37;
ROM_MEM[16013] = 8'hB7;
ROM_MEM[16014] = 8'h18;
ROM_MEM[16015] = 8'h3F;
ROM_MEM[16016] = 8'h96;
ROM_MEM[16017] = 8'h80;
ROM_MEM[16018] = 8'h84;
ROM_MEM[16019] = 8'h10;
ROM_MEM[16020] = 8'h26;
ROM_MEM[16021] = 8'h08;
ROM_MEM[16022] = 8'h96;
ROM_MEM[16023] = 8'h80;
ROM_MEM[16024] = 8'h8A;
ROM_MEM[16025] = 8'h08;
ROM_MEM[16026] = 8'h97;
ROM_MEM[16027] = 8'h80;
ROM_MEM[16028] = 8'h20;
ROM_MEM[16029] = 8'h33;
ROM_MEM[16030] = 8'h96;
ROM_MEM[16031] = 8'h80;
ROM_MEM[16032] = 8'h84;
ROM_MEM[16033] = 8'hF7;
ROM_MEM[16034] = 8'h97;
ROM_MEM[16035] = 8'h80;
ROM_MEM[16036] = 8'h86;
ROM_MEM[16037] = 8'h3F;
ROM_MEM[16038] = 8'h97;
ROM_MEM[16039] = 8'h00;
ROM_MEM[16040] = 8'hBD;
ROM_MEM[16041] = 8'h76;
ROM_MEM[16042] = 8'hA7;
ROM_MEM[16043] = 8'hBD;
ROM_MEM[16044] = 8'h7C;
ROM_MEM[16045] = 8'h45;
ROM_MEM[16046] = 8'h96;
ROM_MEM[16047] = 8'h85;
ROM_MEM[16048] = 8'hB6;
ROM_MEM[16049] = 8'h08;
ROM_MEM[16050] = 8'h00;
ROM_MEM[16051] = 8'h86;
ROM_MEM[16052] = 8'h5A;
ROM_MEM[16053] = 8'hB7;
ROM_MEM[16054] = 8'h00;
ROM_MEM[16055] = 8'h00;
ROM_MEM[16056] = 8'h86;
ROM_MEM[16057] = 8'h06;
ROM_MEM[16058] = 8'h97;
ROM_MEM[16059] = 8'h9F;
ROM_MEM[16060] = 8'h97;
ROM_MEM[16061] = 8'h87;
ROM_MEM[16062] = 8'h7E;
ROM_MEM[16063] = 8'h7D;
ROM_MEM[16064] = 8'h47;
ROM_MEM[16065] = 8'h20;
ROM_MEM[16066] = 8'h00;
ROM_MEM[16067] = 8'h28;
ROM_MEM[16068] = 8'h00;
ROM_MEM[16069] = 8'h01;
ROM_MEM[16070] = 8'h10;
ROM_MEM[16071] = 8'h00;
ROM_MEM[16072] = 8'h10;
ROM_MEM[16073] = 8'h80;
ROM_MEM[16074] = 8'h02;
ROM_MEM[16075] = 8'h40;
ROM_MEM[16076] = 8'h00;
ROM_MEM[16077] = 8'h60;
ROM_MEM[16078] = 8'h00;
ROM_MEM[16079] = 8'h80;
ROM_MEM[16080] = 8'h00;
ROM_MEM[16081] = 8'h86;
ROM_MEM[16082] = 8'h00;
ROM_MEM[16083] = 8'hCE;
ROM_MEM[16084] = 8'h7E;
ROM_MEM[16085] = 8'hC1;
ROM_MEM[16086] = 8'hAE;
ROM_MEM[16087] = 8'hC4;
ROM_MEM[16088] = 8'h31;
ROM_MEM[16089] = 8'h01;
ROM_MEM[16090] = 8'h10;
ROM_MEM[16091] = 8'hAF;
ROM_MEM[16092] = 8'h81;
ROM_MEM[16093] = 8'h31;
ROM_MEM[16094] = 8'hA9;
ROM_MEM[16095] = 8'hFF;
ROM_MEM[16096] = 8'h01;
ROM_MEM[16097] = 8'hAC;
ROM_MEM[16098] = 8'h42;
ROM_MEM[16099] = 8'h25;
ROM_MEM[16100] = 8'hF5;
ROM_MEM[16101] = 8'hAE;
ROM_MEM[16102] = 8'hC4;
ROM_MEM[16103] = 8'h31;
ROM_MEM[16104] = 8'h01;
ROM_MEM[16105] = 8'h10;
ROM_MEM[16106] = 8'hAC;
ROM_MEM[16107] = 8'h81;
ROM_MEM[16108] = 8'h27;
ROM_MEM[16109] = 8'h02;
ROM_MEM[16110] = 8'hAA;
ROM_MEM[16111] = 8'h44;
ROM_MEM[16112] = 8'h31;
ROM_MEM[16113] = 8'hA9;
ROM_MEM[16114] = 8'hFF;
ROM_MEM[16115] = 8'h01;
ROM_MEM[16116] = 8'hAC;
ROM_MEM[16117] = 8'h42;
ROM_MEM[16118] = 8'h25;
ROM_MEM[16119] = 8'hF1;
ROM_MEM[16120] = 8'h33;
ROM_MEM[16121] = 8'h45;
ROM_MEM[16122] = 8'h11;
ROM_MEM[16123] = 8'h83;
ROM_MEM[16124] = 8'h7E;
ROM_MEM[16125] = 8'hCB;
ROM_MEM[16126] = 8'h25;
ROM_MEM[16127] = 8'hD6;
ROM_MEM[16128] = 8'h1F;
ROM_MEM[16129] = 8'h02;
ROM_MEM[16130] = 8'hCE;
ROM_MEM[16131] = 8'h7E;
ROM_MEM[16132] = 8'hCB;
ROM_MEM[16133] = 8'hAE;
ROM_MEM[16134] = 8'hC1;
ROM_MEM[16135] = 8'h1F;
ROM_MEM[16136] = 8'h10;
ROM_MEM[16137] = 8'hE3;
ROM_MEM[16138] = 8'h81;
ROM_MEM[16139] = 8'hAC;
ROM_MEM[16140] = 8'hC4;
ROM_MEM[16141] = 8'h25;
ROM_MEM[16142] = 8'hFA;
ROM_MEM[16143] = 8'hED;
ROM_MEM[16144] = 8'h84;
ROM_MEM[16145] = 8'h27;
ROM_MEM[16146] = 8'h0F;
ROM_MEM[16147] = 8'h1F;
ROM_MEM[16148] = 8'h20;
ROM_MEM[16149] = 8'h8C;
ROM_MEM[16150] = 8'h60;
ROM_MEM[16151] = 8'h10;
ROM_MEM[16152] = 8'h24;
ROM_MEM[16153] = 8'h04;
ROM_MEM[16154] = 8'h8A;
ROM_MEM[16155] = 8'h04;
ROM_MEM[16156] = 8'h20;
ROM_MEM[16157] = 8'h02;
ROM_MEM[16158] = 8'h8A;
ROM_MEM[16159] = 8'h08;
ROM_MEM[16160] = 8'h1F;
ROM_MEM[16161] = 8'h02;
ROM_MEM[16162] = 8'h11;
ROM_MEM[16163] = 8'h83;
ROM_MEM[16164] = 8'h7E;
ROM_MEM[16165] = 8'hCF;
ROM_MEM[16166] = 8'h25;
ROM_MEM[16167] = 8'hDD;
ROM_MEM[16168] = 8'h1F;
ROM_MEM[16169] = 8'h20;
ROM_MEM[16170] = 8'hC6;
ROM_MEM[16171] = 8'h03;
ROM_MEM[16172] = 8'h44;
ROM_MEM[16173] = 8'h24;
ROM_MEM[16174] = 8'h08;
ROM_MEM[16175] = 8'hCE;
ROM_MEM[16176] = 8'hCF;
ROM_MEM[16177] = 8'hA8;
ROM_MEM[16178] = 8'hFF;
ROM_MEM[16179] = 8'h18;
ROM_MEM[16180] = 8'h00;
ROM_MEM[16181] = 8'h20;
ROM_MEM[16182] = 8'h06;
ROM_MEM[16183] = 8'hCE;
ROM_MEM[16184] = 8'h20;
ROM_MEM[16185] = 8'hA8;
ROM_MEM[16186] = 8'hFF;
ROM_MEM[16187] = 8'h18;
ROM_MEM[16188] = 8'h0A;
ROM_MEM[16189] = 8'h8E;
ROM_MEM[16190] = 8'h80;
ROM_MEM[16191] = 8'h00;
ROM_MEM[16192] = 8'h30;
ROM_MEM[16193] = 8'h1F;
ROM_MEM[16194] = 8'h26;
ROM_MEM[16195] = 8'hFC;
ROM_MEM[16196] = 8'hCE;
ROM_MEM[16197] = 8'h00;
ROM_MEM[16198] = 8'h00;
ROM_MEM[16199] = 8'hFF;
ROM_MEM[16200] = 8'h18;
ROM_MEM[16201] = 8'h00;
ROM_MEM[16202] = 8'hFF;
ROM_MEM[16203] = 8'h18;
ROM_MEM[16204] = 8'h0A;
ROM_MEM[16205] = 8'h8E;
ROM_MEM[16206] = 8'h80;
ROM_MEM[16207] = 8'h00;
ROM_MEM[16208] = 8'h5D;
ROM_MEM[16209] = 8'h26;
ROM_MEM[16210] = 8'h04;
ROM_MEM[16211] = 8'h30;
ROM_MEM[16212] = 8'h89;
ROM_MEM[16213] = 8'h7F;
ROM_MEM[16214] = 8'hFF;
ROM_MEM[16215] = 8'h30;
ROM_MEM[16216] = 8'h1F;
ROM_MEM[16217] = 8'h26;
ROM_MEM[16218] = 8'hFC;
ROM_MEM[16219] = 8'h5A;
ROM_MEM[16220] = 8'h2A;
ROM_MEM[16221] = 8'hCE;
ROM_MEM[16222] = 8'h7E;
ROM_MEM[16223] = 8'h7D;
ROM_MEM[16224] = 8'h44;
ROM_MEM[16225] = 8'h7D;
ROM_MEM[16226] = 8'h44;
ROM_MEM[16227] = 8'h74;
ROM_MEM[16228] = 8'h3C;
ROM_MEM[16229] = 8'h76;
ROM_MEM[16230] = 8'h86;
ROM_MEM[16231] = 8'h7B;
ROM_MEM[16232] = 8'hAB;
ROM_MEM[16233] = 8'h7C;
ROM_MEM[16234] = 8'h0D;
ROM_MEM[16235] = 8'h7B;
ROM_MEM[16236] = 8'hBA;
ROM_MEM[16237] = 8'h7B;
ROM_MEM[16238] = 8'hB3;
ROM_MEM[16239] = 8'h7C;
ROM_MEM[16240] = 8'h14;
ROM_MEM[16241] = 8'h7B;
ROM_MEM[16242] = 8'hC2;
ROM_MEM[16243] = 8'h7B;
ROM_MEM[16244] = 8'hDB;
ROM_MEM[16245] = 8'h7C;
ROM_MEM[16246] = 8'h1B;
ROM_MEM[16247] = 8'h7B;
ROM_MEM[16248] = 8'h7E;
ROM_MEM[16249] = 8'h7B;
ROM_MEM[16250] = 8'hFF;
ROM_MEM[16251] = 8'h7B;
ROM_MEM[16252] = 8'hE3;
ROM_MEM[16253] = 8'h7B;
ROM_MEM[16254] = 8'hD4;
ROM_MEM[16255] = 8'h7B;
ROM_MEM[16256] = 8'h6D;
ROM_MEM[16257] = 8'h7B;
ROM_MEM[16258] = 8'h65;
ROM_MEM[16259] = 8'h7B;
ROM_MEM[16260] = 8'hA3;
ROM_MEM[16261] = 8'h7B;
ROM_MEM[16262] = 8'hF1;
ROM_MEM[16263] = 8'h7C;
ROM_MEM[16264] = 8'h06;
ROM_MEM[16265] = 8'h7C;
ROM_MEM[16266] = 8'h40;
ROM_MEM[16267] = 8'h7B;
ROM_MEM[16268] = 8'hCB;
ROM_MEM[16269] = 8'h7B;
ROM_MEM[16270] = 8'h90;
ROM_MEM[16271] = 8'h7B;
ROM_MEM[16272] = 8'h76;
ROM_MEM[16273] = 8'h7B;
ROM_MEM[16274] = 8'hF8;
ROM_MEM[16275] = 8'h7B;
ROM_MEM[16276] = 8'h88;
ROM_MEM[16277] = 8'h7B;
ROM_MEM[16278] = 8'h9A;
ROM_MEM[16279] = 8'h75;
ROM_MEM[16280] = 8'h3C;
ROM_MEM[16281] = 8'h75;
ROM_MEM[16282] = 8'h5D;
ROM_MEM[16283] = 8'h76;
ROM_MEM[16284] = 8'h65;
ROM_MEM[16285] = 8'h76;
ROM_MEM[16286] = 8'h44;
ROM_MEM[16287] = 8'h75;
ROM_MEM[16288] = 8'h7E;
ROM_MEM[16289] = 8'h76;
ROM_MEM[16290] = 8'h02;
ROM_MEM[16291] = 8'h75;
ROM_MEM[16292] = 8'h9F;
ROM_MEM[16293] = 8'h75;
ROM_MEM[16294] = 8'hC0;
ROM_MEM[16295] = 8'h75;
ROM_MEM[16296] = 8'h1B;
ROM_MEM[16297] = 8'h75;
ROM_MEM[16298] = 8'hE1;
ROM_MEM[16299] = 8'h76;
ROM_MEM[16300] = 8'h23;
ROM_MEM[16301] = 8'h74;
ROM_MEM[16302] = 8'h01;
ROM_MEM[16303] = 8'h73;
ROM_MEM[16304] = 8'hF5;
ROM_MEM[16305] = 8'h74;
ROM_MEM[16306] = 8'h0D;
ROM_MEM[16307] = 8'h74;
ROM_MEM[16308] = 8'h35;
ROM_MEM[16309] = 8'h73;
ROM_MEM[16310] = 8'hC5;
ROM_MEM[16311] = 8'h73;
ROM_MEM[16312] = 8'hCB;
ROM_MEM[16313] = 8'h73;
ROM_MEM[16314] = 8'hD7;
ROM_MEM[16315] = 8'h74;
ROM_MEM[16316] = 8'h19;
ROM_MEM[16317] = 8'h73;
ROM_MEM[16318] = 8'hFB;
ROM_MEM[16319] = 8'h74;
ROM_MEM[16320] = 8'h07;
ROM_MEM[16321] = 8'h73;
ROM_MEM[16322] = 8'hB7;
ROM_MEM[16323] = 8'h74;
ROM_MEM[16324] = 8'h20;
ROM_MEM[16325] = 8'h73;
ROM_MEM[16326] = 8'hB0;
ROM_MEM[16327] = 8'h73;
ROM_MEM[16328] = 8'hD1;
ROM_MEM[16329] = 8'h74;
ROM_MEM[16330] = 8'h13;
ROM_MEM[16331] = 8'h73;
ROM_MEM[16332] = 8'hEF;
ROM_MEM[16333] = 8'h73;
ROM_MEM[16334] = 8'hE3;
ROM_MEM[16335] = 8'h73;
ROM_MEM[16336] = 8'hE9;
ROM_MEM[16337] = 8'h74;
ROM_MEM[16338] = 8'h27;
ROM_MEM[16339] = 8'h73;
ROM_MEM[16340] = 8'hDD;
ROM_MEM[16341] = 8'h73;
ROM_MEM[16342] = 8'hBE;
ROM_MEM[16343] = 8'h74;
ROM_MEM[16344] = 8'h2E;
ROM_MEM[16345] = 8'hFF;
ROM_MEM[16346] = 8'hFF;
ROM_MEM[16347] = 8'hFF;
ROM_MEM[16348] = 8'h43;
ROM_MEM[16349] = 8'h4F;
ROM_MEM[16350] = 8'h50;
ROM_MEM[16351] = 8'h59;
ROM_MEM[16352] = 8'h52;
ROM_MEM[16353] = 8'h49;
ROM_MEM[16354] = 8'h47;
ROM_MEM[16355] = 8'h48;
ROM_MEM[16356] = 8'h54;
ROM_MEM[16357] = 8'h20;
ROM_MEM[16358] = 8'h31;
ROM_MEM[16359] = 8'h39;
ROM_MEM[16360] = 8'h38;
ROM_MEM[16361] = 8'h33;
ROM_MEM[16362] = 8'h20;
ROM_MEM[16363] = 8'h41;
ROM_MEM[16364] = 8'h54;
ROM_MEM[16365] = 8'h41;
ROM_MEM[16366] = 8'h52;
ROM_MEM[16367] = 8'h49;
ROM_MEM[16368] = 8'h35;
ROM_MEM[16369] = 8'hE9;
ROM_MEM[16370] = 8'h7E;
ROM_MEM[16371] = 8'h27;
ROM_MEM[16372] = 8'h7E;
ROM_MEM[16373] = 8'h27;
ROM_MEM[16374] = 8'h7E;
ROM_MEM[16375] = 8'h27;
ROM_MEM[16376] = 8'h7D;
ROM_MEM[16377] = 8'hF3;
ROM_MEM[16378] = 8'h7E;
ROM_MEM[16379] = 8'h27;
ROM_MEM[16380] = 8'h7E;
ROM_MEM[16381] = 8'h27;
ROM_MEM[16382] = 8'h7D;
ROM_MEM[16383] = 8'h44;
    end
    
    always @(posedge clk) data <= ROM_MEM[address];
    
    
endmodule
