`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.05.2023 21:37:01
// Design Name: 
// Module Name: matrix_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module matrix_rom (
    input               clk_a,    
    input [9:0]         address_a, 
    output [15:0]       q_a
    
);

reg [7:0] memory0_reg [1023:0];
reg [7:0] memory1_reg [1023:0];
reg [7:0] memory2_reg [1023:0];
reg [7:0] memory3_reg [1023:0];

reg [7:0] memory0;
reg [7:0] memory1;
reg [7:0] memory2;
reg [7:0] memory3;

initial begin
memory0_reg[0   ] <= 8'h09;
memory0_reg[1   ] <= 8'h04;
memory0_reg[2   ] <= 8'h02;
memory0_reg[3   ] <= 8'h08;
memory0_reg[4   ] <= 8'h04;
memory0_reg[5   ] <= 8'h02;
memory0_reg[6   ] <= 8'h08;
memory0_reg[7   ] <= 8'h04;
memory0_reg[8   ] <= 8'h02;
memory0_reg[9   ] <= 8'h08;
memory0_reg[10  ] <= 8'h00;
memory0_reg[11  ] <= 8'h05;
memory0_reg[12  ] <= 8'h02;
memory0_reg[13  ] <= 8'h08;
memory0_reg[14  ] <= 8'h02;
memory0_reg[15  ] <= 8'h08;
memory0_reg[16  ] <= 8'h02;
memory0_reg[17  ] <= 8'h00;
memory0_reg[18  ] <= 8'h09;
memory0_reg[19  ] <= 8'h04;
memory0_reg[20  ] <= 8'h02;
memory0_reg[21  ] <= 8'h08;
memory0_reg[22  ] <= 8'h04;
memory0_reg[23  ] <= 8'h02;
memory0_reg[24  ] <= 8'h08;
memory0_reg[25  ] <= 8'h04;
memory0_reg[26  ] <= 8'h02;
memory0_reg[27  ] <= 8'h08;
memory0_reg[28  ] <= 8'h00;
memory0_reg[29  ] <= 8'h05;
memory0_reg[30  ] <= 8'h02;
memory0_reg[31  ] <= 8'h08;
memory0_reg[32  ] <= 8'h02;
memory0_reg[33  ] <= 8'h08;
memory0_reg[34  ] <= 8'h02;
memory0_reg[35  ] <= 8'h00;
memory0_reg[36  ] <= 8'h09;
memory0_reg[37  ] <= 8'h04;
memory0_reg[38  ] <= 8'h02;
memory0_reg[39  ] <= 8'h08;
memory0_reg[40  ] <= 8'h04;
memory0_reg[41  ] <= 8'h02;
memory0_reg[42  ] <= 8'h08;
memory0_reg[43  ] <= 8'h04;
memory0_reg[44  ] <= 8'h02;
memory0_reg[45  ] <= 8'h08;
memory0_reg[46  ] <= 8'h00;
memory0_reg[47  ] <= 8'h05;
memory0_reg[48  ] <= 8'h02;
memory0_reg[49  ] <= 8'h08;
memory0_reg[50  ] <= 8'h02;
memory0_reg[51  ] <= 8'h08;
memory0_reg[52  ] <= 8'h02;
memory0_reg[53  ] <= 8'h00;
memory0_reg[54  ] <= 8'h00;
memory0_reg[55  ] <= 8'h00;
memory0_reg[56  ] <= 8'h09;
memory0_reg[57  ] <= 8'h04;
memory0_reg[58  ] <= 8'h02;
memory0_reg[59  ] <= 8'h08;
memory0_reg[60  ] <= 8'h04;
memory0_reg[61  ] <= 8'h02;
memory0_reg[62  ] <= 8'h08;
memory0_reg[63  ] <= 8'h04;
memory0_reg[64  ] <= 8'h02;
memory0_reg[65  ] <= 8'h08;
memory0_reg[66  ] <= 8'h00;
memory0_reg[67  ] <= 8'h05;
memory0_reg[68  ] <= 8'h02;
memory0_reg[69  ] <= 8'h08;
memory0_reg[70  ] <= 8'h02;
memory0_reg[71  ] <= 8'h08;
memory0_reg[72  ] <= 8'h02;
memory0_reg[73  ] <= 8'h00;
memory0_reg[74  ] <= 8'h09;
memory0_reg[75  ] <= 8'h04;
memory0_reg[76  ] <= 8'h02;
memory0_reg[77  ] <= 8'h08;
memory0_reg[78  ] <= 8'h04;
memory0_reg[79  ] <= 8'h02;
memory0_reg[80  ] <= 8'h08;
memory0_reg[81  ] <= 8'h04;
memory0_reg[82  ] <= 8'h02;
memory0_reg[83  ] <= 8'h08;
memory0_reg[84  ] <= 8'h00;
memory0_reg[85  ] <= 8'h05;
memory0_reg[86  ] <= 8'h02;
memory0_reg[87  ] <= 8'h08;
memory0_reg[88  ] <= 8'h02;
memory0_reg[89  ] <= 8'h08;
memory0_reg[90  ] <= 8'h02;
memory0_reg[91  ] <= 8'h00;
memory0_reg[92  ] <= 8'h09;
memory0_reg[93  ] <= 8'h04;
memory0_reg[94  ] <= 8'h02;
memory0_reg[95  ] <= 8'h08;
memory0_reg[96  ] <= 8'h04;
memory0_reg[97  ] <= 8'h02;
memory0_reg[98  ] <= 8'h08;
memory0_reg[99  ] <= 8'h04;
memory0_reg[100 ] <= 8'h02;
memory0_reg[101 ] <= 8'h08;
memory0_reg[102 ] <= 8'h00;
memory0_reg[103 ] <= 8'h05;
memory0_reg[104 ] <= 8'h02;
memory0_reg[105 ] <= 8'h08;
memory0_reg[106 ] <= 8'h02;
memory0_reg[107 ] <= 8'h08;
memory0_reg[108 ] <= 8'h02;
memory0_reg[109 ] <= 8'h00;
memory0_reg[110 ] <= 8'h00;
memory0_reg[111 ] <= 8'h00;
memory0_reg[112 ] <= 8'h09;
memory0_reg[113 ] <= 8'h04;
memory0_reg[114 ] <= 8'h02;
memory0_reg[115 ] <= 8'h08;
memory0_reg[116 ] <= 8'h04;
memory0_reg[117 ] <= 8'h02;
memory0_reg[118 ] <= 8'h08;
memory0_reg[119 ] <= 8'h04;
memory0_reg[120 ] <= 8'h02;
memory0_reg[121 ] <= 8'h08;
memory0_reg[122 ] <= 8'h00;
memory0_reg[123 ] <= 8'h05;
memory0_reg[124 ] <= 8'h02;
memory0_reg[125 ] <= 8'h08;
memory0_reg[126 ] <= 8'h02;
memory0_reg[127 ] <= 8'h08;
memory0_reg[128 ] <= 8'h02;
memory0_reg[129 ] <= 8'h00;
memory0_reg[130 ] <= 8'h09;
memory0_reg[131 ] <= 8'h04;
memory0_reg[132 ] <= 8'h02;
memory0_reg[133 ] <= 8'h08;
memory0_reg[134 ] <= 8'h04;
memory0_reg[135 ] <= 8'h02;
memory0_reg[136 ] <= 8'h08;
memory0_reg[137 ] <= 8'h04;
memory0_reg[138 ] <= 8'h02;
memory0_reg[139 ] <= 8'h08;
memory0_reg[140 ] <= 8'h00;
memory0_reg[141 ] <= 8'h05;
memory0_reg[142 ] <= 8'h02;
memory0_reg[143 ] <= 8'h08;
memory0_reg[144 ] <= 8'h02;
memory0_reg[145 ] <= 8'h08;
memory0_reg[146 ] <= 8'h02;
memory0_reg[147 ] <= 8'h00;
memory0_reg[148 ] <= 8'h09;
memory0_reg[149 ] <= 8'h04;
memory0_reg[150 ] <= 8'h02;
memory0_reg[151 ] <= 8'h08;
memory0_reg[152 ] <= 8'h04;
memory0_reg[153 ] <= 8'h02;
memory0_reg[154 ] <= 8'h08;
memory0_reg[155 ] <= 8'h04;
memory0_reg[156 ] <= 8'h02;
memory0_reg[157 ] <= 8'h08;
memory0_reg[158 ] <= 8'h00;
memory0_reg[159 ] <= 8'h05;
memory0_reg[160 ] <= 8'h02;
memory0_reg[161 ] <= 8'h08;
memory0_reg[162 ] <= 8'h02;
memory0_reg[163 ] <= 8'h08;
memory0_reg[164 ] <= 8'h02;
memory0_reg[165 ] <= 8'h00;
memory0_reg[166 ] <= 8'h00;
memory0_reg[167 ] <= 8'h00;
memory0_reg[168 ] <= 8'h09;
memory0_reg[169 ] <= 8'h04;
memory0_reg[170 ] <= 8'h02;
memory0_reg[171 ] <= 8'h08;
memory0_reg[172 ] <= 8'h04;
memory0_reg[173 ] <= 8'h02;
memory0_reg[174 ] <= 8'h08;
memory0_reg[175 ] <= 8'h04;
memory0_reg[176 ] <= 8'h02;
memory0_reg[177 ] <= 8'h00;
memory0_reg[178 ] <= 8'h09;
memory0_reg[179 ] <= 8'h04;
memory0_reg[180 ] <= 8'h02;
memory0_reg[181 ] <= 8'h08;
memory0_reg[182 ] <= 8'h04;
memory0_reg[183 ] <= 8'h02;
memory0_reg[184 ] <= 8'h08;
memory0_reg[185 ] <= 8'h04;
memory0_reg[186 ] <= 8'h02;
memory0_reg[187 ] <= 8'h00;
memory0_reg[188 ] <= 8'h09;
memory0_reg[189 ] <= 8'h04;
memory0_reg[190 ] <= 8'h02;
memory0_reg[191 ] <= 8'h08;
memory0_reg[192 ] <= 8'h04;
memory0_reg[193 ] <= 8'h02;
memory0_reg[194 ] <= 8'h08;
memory0_reg[195 ] <= 8'h04;
memory0_reg[196 ] <= 8'h02;
memory0_reg[197 ] <= 8'h00;
memory0_reg[198 ] <= 8'h00;
memory0_reg[199 ] <= 8'h00;
memory0_reg[200 ] <= 8'h00;
memory0_reg[201 ] <= 8'h00;
memory0_reg[202 ] <= 8'h00;
memory0_reg[203 ] <= 8'h00;
memory0_reg[204 ] <= 8'h00;
memory0_reg[205 ] <= 8'h00;
memory0_reg[206 ] <= 8'h00;
memory0_reg[207 ] <= 8'h00;
memory0_reg[208 ] <= 8'h00;
memory0_reg[209 ] <= 8'h00;
memory0_reg[210 ] <= 8'h00;
memory0_reg[211 ] <= 8'h00;
memory0_reg[212 ] <= 8'h00;
memory0_reg[213 ] <= 8'h00;
memory0_reg[214 ] <= 8'h00;
memory0_reg[215 ] <= 8'h00;
memory0_reg[216 ] <= 8'h00;
memory0_reg[217 ] <= 8'h00;
memory0_reg[218 ] <= 8'h00;
memory0_reg[219 ] <= 8'h00;
memory0_reg[220 ] <= 8'h00;
memory0_reg[221 ] <= 8'h00;
memory0_reg[222 ] <= 8'h00;
memory0_reg[223 ] <= 8'h00;
memory0_reg[224 ] <= 8'h00;
memory0_reg[225 ] <= 8'h00;
memory0_reg[226 ] <= 8'h00;
memory0_reg[227 ] <= 8'h00;
memory0_reg[228 ] <= 8'h00;
memory0_reg[229 ] <= 8'h00;
memory0_reg[230 ] <= 8'h00;
memory0_reg[231 ] <= 8'h00;
memory0_reg[232 ] <= 8'h00;
memory0_reg[233 ] <= 8'h00;
memory0_reg[234 ] <= 8'h00;
memory0_reg[235 ] <= 8'h00;
memory0_reg[236 ] <= 8'h00;
memory0_reg[237 ] <= 8'h00;
memory0_reg[238 ] <= 8'h00;
memory0_reg[239 ] <= 8'h00;
memory0_reg[240 ] <= 8'h00;
memory0_reg[241 ] <= 8'h00;
memory0_reg[242 ] <= 8'h00;
memory0_reg[243 ] <= 8'h00;
memory0_reg[244 ] <= 8'h00;
memory0_reg[245 ] <= 8'h00;
memory0_reg[246 ] <= 8'h00;
memory0_reg[247 ] <= 8'h00;
memory0_reg[248 ] <= 8'h00;
memory0_reg[249 ] <= 8'h00;
memory0_reg[250 ] <= 8'h00;
memory0_reg[251 ] <= 8'h00;
memory0_reg[252 ] <= 8'h00;
memory0_reg[253 ] <= 8'h00;
memory0_reg[254 ] <= 8'h00;
memory0_reg[255 ] <= 8'h00;
memory0_reg[256 ] <= 8'h04;
memory0_reg[257 ] <= 8'h09;
memory0_reg[258 ] <= 8'h02;
memory0_reg[259 ] <= 8'h08;
memory0_reg[260 ] <= 8'h02;
memory0_reg[261 ] <= 8'h08;
memory0_reg[262 ] <= 8'h02;
memory0_reg[263 ] <= 8'h00;
memory0_reg[264 ] <= 8'h09;
memory0_reg[265 ] <= 8'h02;
memory0_reg[266 ] <= 8'h08;
memory0_reg[267 ] <= 8'h02;
memory0_reg[268 ] <= 8'h08;
memory0_reg[269 ] <= 8'h02;
memory0_reg[270 ] <= 8'h00;
memory0_reg[271 ] <= 8'h09;
memory0_reg[272 ] <= 8'h02;
memory0_reg[273 ] <= 8'h08;
memory0_reg[274 ] <= 8'h02;
memory0_reg[275 ] <= 8'h08;
memory0_reg[276 ] <= 8'h02;
memory0_reg[277 ] <= 8'h00;
memory0_reg[278 ] <= 8'h09;
memory0_reg[279 ] <= 8'h02;
memory0_reg[280 ] <= 8'h08;
memory0_reg[281 ] <= 8'h02;
memory0_reg[282 ] <= 8'h08;
memory0_reg[283 ] <= 8'h02;
memory0_reg[284 ] <= 8'h00;
memory0_reg[285 ] <= 8'h09;
memory0_reg[286 ] <= 8'h02;
memory0_reg[287 ] <= 8'h08;
memory0_reg[288 ] <= 8'h02;
memory0_reg[289 ] <= 8'h08;
memory0_reg[290 ] <= 8'h02;
memory0_reg[291 ] <= 8'h00;
memory0_reg[292 ] <= 8'h09;
memory0_reg[293 ] <= 8'h02;
memory0_reg[294 ] <= 8'h08;
memory0_reg[295 ] <= 8'h02;
memory0_reg[296 ] <= 8'h08;
memory0_reg[297 ] <= 8'h02;
memory0_reg[298 ] <= 8'h00;
memory0_reg[299 ] <= 8'h09;
memory0_reg[300 ] <= 8'h02;
memory0_reg[301 ] <= 8'h08;
memory0_reg[302 ] <= 8'h02;
memory0_reg[303 ] <= 8'h08;
memory0_reg[304 ] <= 8'h02;
memory0_reg[305 ] <= 8'h00;
memory0_reg[306 ] <= 8'h09;
memory0_reg[307 ] <= 8'h02;
memory0_reg[308 ] <= 8'h08;
memory0_reg[309 ] <= 8'h02;
memory0_reg[310 ] <= 8'h08;
memory0_reg[311 ] <= 8'h02;
memory0_reg[312 ] <= 8'h00;
memory0_reg[313 ] <= 8'h09;
memory0_reg[314 ] <= 8'h02;
memory0_reg[315 ] <= 8'h08;
memory0_reg[316 ] <= 8'h02;
memory0_reg[317 ] <= 8'h08;
memory0_reg[318 ] <= 8'h02;
memory0_reg[319 ] <= 8'h00;
memory0_reg[320 ] <= 8'h04;
memory0_reg[321 ] <= 8'h00;
memory0_reg[322 ] <= 8'h08;
memory0_reg[323 ] <= 8'h02;
memory0_reg[324 ] <= 8'h08;
memory0_reg[325 ] <= 8'h02;
memory0_reg[326 ] <= 8'h08;
memory0_reg[327 ] <= 8'h02;
memory0_reg[328 ] <= 8'h00;
memory0_reg[329 ] <= 8'h00;
memory0_reg[330 ] <= 8'h08;
memory0_reg[331 ] <= 8'h02;
memory0_reg[332 ] <= 8'h08;
memory0_reg[333 ] <= 8'h02;
memory0_reg[334 ] <= 8'h08;
memory0_reg[335 ] <= 8'h02;
memory0_reg[336 ] <= 8'h00;
memory0_reg[337 ] <= 8'h00;
memory0_reg[338 ] <= 8'h08;
memory0_reg[339 ] <= 8'h02;
memory0_reg[340 ] <= 8'h08;
memory0_reg[341 ] <= 8'h02;
memory0_reg[342 ] <= 8'h08;
memory0_reg[343 ] <= 8'h02;
memory0_reg[344 ] <= 8'h00;
memory0_reg[345 ] <= 8'h09;
memory0_reg[346 ] <= 8'h02;
memory0_reg[347 ] <= 8'h00;
memory0_reg[348 ] <= 8'h08;
memory0_reg[349 ] <= 8'h00;
memory0_reg[350 ] <= 8'h00;
memory0_reg[351 ] <= 8'h00;
memory0_reg[352 ] <= 8'h04;
memory0_reg[353 ] <= 8'h00;
memory0_reg[354 ] <= 8'h00;
memory0_reg[355 ] <= 8'h00;
memory0_reg[356 ] <= 8'h02;
memory0_reg[357 ] <= 8'h00;
memory0_reg[358 ] <= 8'h00;
memory0_reg[359 ] <= 8'h00;
memory0_reg[360 ] <= 8'h01;
memory0_reg[361 ] <= 8'h00;
memory0_reg[362 ] <= 8'h00;
memory0_reg[363 ] <= 8'h00;
memory0_reg[364 ] <= 8'h00;
memory0_reg[365 ] <= 8'h00;
memory0_reg[366 ] <= 8'h00;
memory0_reg[367 ] <= 8'h00;
memory0_reg[368 ] <= 8'h00;
memory0_reg[369 ] <= 8'h00;
memory0_reg[370 ] <= 8'h00;
memory0_reg[371 ] <= 8'h00;
memory0_reg[372 ] <= 8'h09;
memory0_reg[373 ] <= 8'h04;
memory0_reg[374 ] <= 8'h02;
memory0_reg[375 ] <= 8'h00;
memory0_reg[376 ] <= 8'h08;
memory0_reg[377 ] <= 8'h04;
memory0_reg[378 ] <= 8'h02;
memory0_reg[379 ] <= 8'h00;
memory0_reg[380 ] <= 8'h09;
memory0_reg[381 ] <= 8'h04;
memory0_reg[382 ] <= 8'h02;
memory0_reg[383 ] <= 8'h00;
memory0_reg[384 ] <= 8'h04;
memory0_reg[385 ] <= 8'h00;
memory0_reg[386 ] <= 8'h08;
memory0_reg[387 ] <= 8'h02;
memory0_reg[388 ] <= 8'h08;
memory0_reg[389 ] <= 8'h02;
memory0_reg[390 ] <= 8'h08;
memory0_reg[391 ] <= 8'h02;
memory0_reg[392 ] <= 8'h00;
memory0_reg[393 ] <= 8'h00;
memory0_reg[394 ] <= 8'h08;
memory0_reg[395 ] <= 8'h02;
memory0_reg[396 ] <= 8'h08;
memory0_reg[397 ] <= 8'h02;
memory0_reg[398 ] <= 8'h08;
memory0_reg[399 ] <= 8'h02;
memory0_reg[400 ] <= 8'h00;
memory0_reg[401 ] <= 8'h00;
memory0_reg[402 ] <= 8'h08;
memory0_reg[403 ] <= 8'h02;
memory0_reg[404 ] <= 8'h08;
memory0_reg[405 ] <= 8'h02;
memory0_reg[406 ] <= 8'h08;
memory0_reg[407 ] <= 8'h02;
memory0_reg[408 ] <= 8'h00;
memory0_reg[409 ] <= 8'h00;
memory0_reg[410 ] <= 8'h00;
memory0_reg[411 ] <= 8'h00;
memory0_reg[412 ] <= 8'h09;
memory0_reg[413 ] <= 8'h04;
memory0_reg[414 ] <= 8'h02;
memory0_reg[415 ] <= 8'h00;
memory0_reg[416 ] <= 8'h08;
memory0_reg[417 ] <= 8'h04;
memory0_reg[418 ] <= 8'h02;
memory0_reg[419 ] <= 8'h00;
memory0_reg[420 ] <= 8'h09;
memory0_reg[421 ] <= 8'h04;
memory0_reg[422 ] <= 8'h02;
memory0_reg[423 ] <= 8'h00;
memory0_reg[424 ] <= 8'h08;
memory0_reg[425 ] <= 8'h04;
memory0_reg[426 ] <= 8'h02;
memory0_reg[427 ] <= 8'h00;
memory0_reg[428 ] <= 8'h09;
memory0_reg[429 ] <= 8'h04;
memory0_reg[430 ] <= 8'h02;
memory0_reg[431 ] <= 8'h00;
memory0_reg[432 ] <= 8'h08;
memory0_reg[433 ] <= 8'h04;
memory0_reg[434 ] <= 8'h02;
memory0_reg[435 ] <= 8'h00;
memory0_reg[436 ] <= 8'h04;
memory0_reg[437 ] <= 8'h09;
memory0_reg[438 ] <= 8'h02;
memory0_reg[439 ] <= 8'h08;
memory0_reg[440 ] <= 8'h02;
memory0_reg[441 ] <= 8'h08;
memory0_reg[442 ] <= 8'h02;
memory0_reg[443 ] <= 8'h00;
memory0_reg[444 ] <= 8'h09;
memory0_reg[445 ] <= 8'h02;
memory0_reg[446 ] <= 8'h08;
memory0_reg[447 ] <= 8'h02;
memory0_reg[448 ] <= 8'h08;
memory0_reg[449 ] <= 8'h02;
memory0_reg[450 ] <= 8'h00;
memory0_reg[451 ] <= 8'h09;
memory0_reg[452 ] <= 8'h02;
memory0_reg[453 ] <= 8'h08;
memory0_reg[454 ] <= 8'h02;
memory0_reg[455 ] <= 8'h08;
memory0_reg[456 ] <= 8'h02;
memory0_reg[457 ] <= 8'h00;
memory0_reg[458 ] <= 8'h09;
memory0_reg[459 ] <= 8'h02;
memory0_reg[460 ] <= 8'h00;
memory0_reg[461 ] <= 8'h09;
memory0_reg[462 ] <= 8'h02;
memory0_reg[463 ] <= 8'h00;
memory0_reg[464 ] <= 8'h09;
memory0_reg[465 ] <= 8'h02;
memory0_reg[466 ] <= 8'h00;
memory0_reg[467 ] <= 8'h09;
memory0_reg[468 ] <= 8'h02;
memory0_reg[469 ] <= 8'h00;
memory0_reg[470 ] <= 8'h09;
memory0_reg[471 ] <= 8'h02;
memory0_reg[472 ] <= 8'h00;
memory0_reg[473 ] <= 8'h00;
memory0_reg[474 ] <= 8'h00;
memory0_reg[475 ] <= 8'h00;
memory0_reg[476 ] <= 8'h00;
memory0_reg[477 ] <= 8'h00;
memory0_reg[478 ] <= 8'h00;
memory0_reg[479 ] <= 8'h00;
memory0_reg[480 ] <= 8'h00;
memory0_reg[481 ] <= 8'h00;
memory0_reg[482 ] <= 8'h00;
memory0_reg[483 ] <= 8'h00;
memory0_reg[484 ] <= 8'h00;
memory0_reg[485 ] <= 8'h00;
memory0_reg[486 ] <= 8'h00;
memory0_reg[487 ] <= 8'h00;
memory0_reg[488 ] <= 8'h00;
memory0_reg[489 ] <= 8'h00;
memory0_reg[490 ] <= 8'h00;
memory0_reg[491 ] <= 8'h00;
memory0_reg[492 ] <= 8'h00;
memory0_reg[493 ] <= 8'h00;
memory0_reg[494 ] <= 8'h00;
memory0_reg[495 ] <= 8'h00;
memory0_reg[496 ] <= 8'h00;
memory0_reg[497 ] <= 8'h00;
memory0_reg[498 ] <= 8'h00;
memory0_reg[499 ] <= 8'h00;
memory0_reg[500 ] <= 8'h00;
memory0_reg[501 ] <= 8'h00;
memory0_reg[502 ] <= 8'h00;
memory0_reg[503 ] <= 8'h00;
memory0_reg[504 ] <= 8'h00;
memory0_reg[505 ] <= 8'h00;
memory0_reg[506 ] <= 8'h00;
memory0_reg[507 ] <= 8'h00;
memory0_reg[508 ] <= 8'h00;
memory0_reg[509 ] <= 8'h00;
memory0_reg[510 ] <= 8'h00;
memory0_reg[511 ] <= 8'h00;
memory0_reg[512 ] <= 8'h00;
memory0_reg[513 ] <= 8'h00;
memory0_reg[514 ] <= 8'h00;
memory0_reg[515 ] <= 8'h00;
memory0_reg[516 ] <= 8'h00;
memory0_reg[517 ] <= 8'h00;
memory0_reg[518 ] <= 8'h00;
memory0_reg[519 ] <= 8'h00;
memory0_reg[520 ] <= 8'h00;
memory0_reg[521 ] <= 8'h00;
memory0_reg[522 ] <= 8'h00;
memory0_reg[523 ] <= 8'h00;
memory0_reg[524 ] <= 8'h00;
memory0_reg[525 ] <= 8'h00;
memory0_reg[526 ] <= 8'h00;
memory0_reg[527 ] <= 8'h00;
memory0_reg[528 ] <= 8'h00;
memory0_reg[529 ] <= 8'h00;
memory0_reg[530 ] <= 8'h00;
memory0_reg[531 ] <= 8'h00;
memory0_reg[532 ] <= 8'h00;
memory0_reg[533 ] <= 8'h00;
memory0_reg[534 ] <= 8'h00;
memory0_reg[535 ] <= 8'h00;
memory0_reg[536 ] <= 8'h04;
memory0_reg[537 ] <= 8'h09;
memory0_reg[538 ] <= 8'h02;
memory0_reg[539 ] <= 8'h00;
memory0_reg[540 ] <= 8'h09;
memory0_reg[541 ] <= 8'h02;
memory0_reg[542 ] <= 8'h00;
memory0_reg[543 ] <= 8'h00;
memory0_reg[544 ] <= 8'h04;
memory0_reg[545 ] <= 8'h09;
memory0_reg[546 ] <= 8'h02;
memory0_reg[547 ] <= 8'h08;
memory0_reg[548 ] <= 8'h02;
memory0_reg[549 ] <= 8'h00;
memory0_reg[550 ] <= 8'h00;
memory0_reg[551 ] <= 8'h00;
memory0_reg[552 ] <= 8'h09;
memory0_reg[553 ] <= 8'h02;
memory0_reg[554 ] <= 8'h00;
memory0_reg[555 ] <= 8'h09;
memory0_reg[556 ] <= 8'h02;
memory0_reg[557 ] <= 8'h00;
memory0_reg[558 ] <= 8'h09;
memory0_reg[559 ] <= 8'h02;
memory0_reg[560 ] <= 8'h00;
memory0_reg[561 ] <= 8'h09;
memory0_reg[562 ] <= 8'h04;
memory0_reg[563 ] <= 8'h02;
memory0_reg[564 ] <= 8'h04;
memory0_reg[565 ] <= 8'h08;
memory0_reg[566 ] <= 8'h02;
memory0_reg[567 ] <= 8'h08;
memory0_reg[568 ] <= 8'h02;
memory0_reg[569 ] <= 8'h00;
memory0_reg[570 ] <= 8'h09;
memory0_reg[571 ] <= 8'h04;
memory0_reg[572 ] <= 8'h02;
memory0_reg[573 ] <= 8'h04;
memory0_reg[574 ] <= 8'h08;
memory0_reg[575 ] <= 8'h02;
memory0_reg[576 ] <= 8'h08;
memory0_reg[577 ] <= 8'h02;
memory0_reg[578 ] <= 8'h00;
memory0_reg[579 ] <= 8'h09;
memory0_reg[580 ] <= 8'h02;
memory0_reg[581 ] <= 8'h08;
memory0_reg[582 ] <= 8'h02;
memory0_reg[583 ] <= 8'h08;
memory0_reg[584 ] <= 8'h04;
memory0_reg[585 ] <= 8'h02;
memory0_reg[586 ] <= 8'h00;
memory0_reg[587 ] <= 8'h04;
memory0_reg[588 ] <= 8'h09;
memory0_reg[589 ] <= 8'h02;
memory0_reg[590 ] <= 8'h08;
memory0_reg[591 ] <= 8'h02;
memory0_reg[592 ] <= 8'h08;
memory0_reg[593 ] <= 8'h04;
memory0_reg[594 ] <= 8'h02;
memory0_reg[595 ] <= 8'h00;
memory0_reg[596 ] <= 8'h04;
memory0_reg[597 ] <= 8'h09;
memory0_reg[598 ] <= 8'h02;
memory0_reg[599 ] <= 8'h00;
memory0_reg[600 ] <= 8'h08;
memory0_reg[601 ] <= 8'h05;
memory0_reg[602 ] <= 8'h02;
memory0_reg[603 ] <= 8'h04;
memory0_reg[604 ] <= 8'h02;
memory0_reg[605 ] <= 8'h04;
memory0_reg[606 ] <= 8'h02;
memory0_reg[607 ] <= 8'h00;
memory0_reg[608 ] <= 8'h09;
memory0_reg[609 ] <= 8'h02;
memory0_reg[610 ] <= 8'h08;
memory0_reg[611 ] <= 8'h02;
memory0_reg[612 ] <= 8'h08;
memory0_reg[613 ] <= 8'h02;
memory0_reg[614 ] <= 8'h00;
memory0_reg[615 ] <= 8'h09;
memory0_reg[616 ] <= 8'h02;
memory0_reg[617 ] <= 8'h08;
memory0_reg[618 ] <= 8'h02;
memory0_reg[619 ] <= 8'h08;
memory0_reg[620 ] <= 8'h02;
memory0_reg[621 ] <= 8'h00;
memory0_reg[622 ] <= 8'h00;
memory0_reg[623 ] <= 8'h08;
memory0_reg[624 ] <= 8'h02;
memory0_reg[625 ] <= 8'h08;
memory0_reg[626 ] <= 8'h02;
memory0_reg[627 ] <= 8'h08;
memory0_reg[628 ] <= 8'h02;
memory0_reg[629 ] <= 8'h00;
memory0_reg[630 ] <= 8'h00;
memory0_reg[631 ] <= 8'h00;
memory0_reg[632 ] <= 8'h04;
memory0_reg[633 ] <= 8'h09;
memory0_reg[634 ] <= 8'h02;
memory0_reg[635 ] <= 8'h00;
memory0_reg[636 ] <= 8'h09;
memory0_reg[637 ] <= 8'h02;
memory0_reg[638 ] <= 8'h08;
memory0_reg[639 ] <= 8'h02;
memory0_reg[640 ] <= 8'h00;
memory0_reg[641 ] <= 8'h09;
memory0_reg[642 ] <= 8'h02;
memory0_reg[643 ] <= 8'h08;
memory0_reg[644 ] <= 8'h02;
memory0_reg[645 ] <= 8'h00;
memory0_reg[646 ] <= 8'h00;
memory0_reg[647 ] <= 8'h08;
memory0_reg[648 ] <= 8'h02;
memory0_reg[649 ] <= 8'h08;
memory0_reg[650 ] <= 8'h02;
memory0_reg[651 ] <= 8'h00;
memory0_reg[652 ] <= 8'h04;
memory0_reg[653 ] <= 8'h09;
memory0_reg[654 ] <= 8'h02;
memory0_reg[655 ] <= 8'h00;
memory0_reg[656 ] <= 8'h08;
memory0_reg[657 ] <= 8'h05;
memory0_reg[658 ] <= 8'h02;
memory0_reg[659 ] <= 8'h04;
memory0_reg[660 ] <= 8'h02;
memory0_reg[661 ] <= 8'h04;
memory0_reg[662 ] <= 8'h02;
memory0_reg[663 ] <= 8'h00;
memory0_reg[664 ] <= 8'h04;
memory0_reg[665 ] <= 8'h09;
memory0_reg[666 ] <= 8'h02;
memory0_reg[667 ] <= 8'h08;
memory0_reg[668 ] <= 8'h02;
memory0_reg[669 ] <= 8'h08;
memory0_reg[670 ] <= 8'h02;
memory0_reg[671 ] <= 8'h00;
memory0_reg[672 ] <= 8'h09;
memory0_reg[673 ] <= 8'h02;
memory0_reg[674 ] <= 8'h08;
memory0_reg[675 ] <= 8'h02;
memory0_reg[676 ] <= 8'h08;
memory0_reg[677 ] <= 8'h02;
memory0_reg[678 ] <= 8'h00;
memory0_reg[679 ] <= 8'h00;
memory0_reg[680 ] <= 8'h08;
memory0_reg[681 ] <= 8'h02;
memory0_reg[682 ] <= 8'h08;
memory0_reg[683 ] <= 8'h02;
memory0_reg[684 ] <= 8'h08;
memory0_reg[685 ] <= 8'h02;
memory0_reg[686 ] <= 8'h00;
memory0_reg[687 ] <= 8'h00;
memory0_reg[688 ] <= 8'h05;
memory0_reg[689 ] <= 8'h08;
memory0_reg[690 ] <= 8'h02;
memory0_reg[691 ] <= 8'h08;
memory0_reg[692 ] <= 8'h02;
memory0_reg[693 ] <= 8'h08;
memory0_reg[694 ] <= 8'h02;
memory0_reg[695 ] <= 8'h00;
memory0_reg[696 ] <= 8'h08;
memory0_reg[697 ] <= 8'h05;
memory0_reg[698 ] <= 8'h02;
memory0_reg[699 ] <= 8'h00;
memory0_reg[700 ] <= 8'h08;
memory0_reg[701 ] <= 8'h05;
memory0_reg[702 ] <= 8'h02;
memory0_reg[703 ] <= 8'h00;
memory0_reg[704 ] <= 8'h08;
memory0_reg[705 ] <= 8'h05;
memory0_reg[706 ] <= 8'h02;
memory0_reg[707 ] <= 8'h00;
memory0_reg[708 ] <= 8'h00;
memory0_reg[709 ] <= 8'h00;
memory0_reg[710 ] <= 8'h00;
memory0_reg[711 ] <= 8'h00;
memory0_reg[712 ] <= 8'h00;
memory0_reg[713 ] <= 8'h00;
memory0_reg[714 ] <= 8'h00;
memory0_reg[715 ] <= 8'h00;
memory0_reg[716 ] <= 8'h00;
memory0_reg[717 ] <= 8'h00;
memory0_reg[718 ] <= 8'h00;
memory0_reg[719 ] <= 8'h00;
memory0_reg[720 ] <= 8'h00;
memory0_reg[721 ] <= 8'h00;
memory0_reg[722 ] <= 8'h00;
memory0_reg[723 ] <= 8'h00;
memory0_reg[724 ] <= 8'h00;
memory0_reg[725 ] <= 8'h00;
memory0_reg[726 ] <= 8'h00;
memory0_reg[727 ] <= 8'h00;
memory0_reg[728 ] <= 8'h00;
memory0_reg[729 ] <= 8'h00;
memory0_reg[730 ] <= 8'h00;
memory0_reg[731 ] <= 8'h00;
memory0_reg[732 ] <= 8'h00;
memory0_reg[733 ] <= 8'h00;
memory0_reg[734 ] <= 8'h00;
memory0_reg[735 ] <= 8'h00;
memory0_reg[736 ] <= 8'h00;
memory0_reg[737 ] <= 8'h00;
memory0_reg[738 ] <= 8'h00;
memory0_reg[739 ] <= 8'h00;
memory0_reg[740 ] <= 8'h00;
memory0_reg[741 ] <= 8'h00;
memory0_reg[742 ] <= 8'h00;
memory0_reg[743 ] <= 8'h00;
memory0_reg[744 ] <= 8'h00;
memory0_reg[745 ] <= 8'h00;
memory0_reg[746 ] <= 8'h00;
memory0_reg[747 ] <= 8'h00;
memory0_reg[748 ] <= 8'h00;
memory0_reg[749 ] <= 8'h00;
memory0_reg[750 ] <= 8'h00;
memory0_reg[751 ] <= 8'h00;
memory0_reg[752 ] <= 8'h00;
memory0_reg[753 ] <= 8'h00;
memory0_reg[754 ] <= 8'h00;
memory0_reg[755 ] <= 8'h00;
memory0_reg[756 ] <= 8'h00;
memory0_reg[757 ] <= 8'h00;
memory0_reg[758 ] <= 8'h00;
memory0_reg[759 ] <= 8'h00;
memory0_reg[760 ] <= 8'h00;
memory0_reg[761 ] <= 8'h00;
memory0_reg[762 ] <= 8'h00;
memory0_reg[763 ] <= 8'h00;
memory0_reg[764 ] <= 8'h00;
memory0_reg[765 ] <= 8'h00;
memory0_reg[766 ] <= 8'h00;
memory0_reg[767 ] <= 8'h00;
memory0_reg[768 ] <= 8'h00;
memory0_reg[769 ] <= 8'h00;
memory0_reg[770 ] <= 8'h00;
memory0_reg[771 ] <= 8'h00;
memory0_reg[772 ] <= 8'h00;
memory0_reg[773 ] <= 8'h00;
memory0_reg[774 ] <= 8'h00;
memory0_reg[775 ] <= 8'h00;
memory0_reg[776 ] <= 8'h00;
memory0_reg[777 ] <= 8'h00;
memory0_reg[778 ] <= 8'h00;
memory0_reg[779 ] <= 8'h00;
memory0_reg[780 ] <= 8'h00;
memory0_reg[781 ] <= 8'h00;
memory0_reg[782 ] <= 8'h00;
memory0_reg[783 ] <= 8'h00;
memory0_reg[784 ] <= 8'h00;
memory0_reg[785 ] <= 8'h00;
memory0_reg[786 ] <= 8'h00;
memory0_reg[787 ] <= 8'h00;
memory0_reg[788 ] <= 8'h00;
memory0_reg[789 ] <= 8'h00;
memory0_reg[790 ] <= 8'h00;
memory0_reg[791 ] <= 8'h00;
memory0_reg[792 ] <= 8'h00;
memory0_reg[793 ] <= 8'h00;
memory0_reg[794 ] <= 8'h00;
memory0_reg[795 ] <= 8'h00;
memory0_reg[796 ] <= 8'h00;
memory0_reg[797 ] <= 8'h00;
memory0_reg[798 ] <= 8'h00;
memory0_reg[799 ] <= 8'h00;
memory0_reg[800 ] <= 8'h00;
memory0_reg[801 ] <= 8'h00;
memory0_reg[802 ] <= 8'h00;
memory0_reg[803 ] <= 8'h00;
memory0_reg[804 ] <= 8'h00;
memory0_reg[805 ] <= 8'h00;
memory0_reg[806 ] <= 8'h00;
memory0_reg[807 ] <= 8'h00;
memory0_reg[808 ] <= 8'h00;
memory0_reg[809 ] <= 8'h00;
memory0_reg[810 ] <= 8'h00;
memory0_reg[811 ] <= 8'h00;
memory0_reg[812 ] <= 8'h00;
memory0_reg[813 ] <= 8'h00;
memory0_reg[814 ] <= 8'h00;
memory0_reg[815 ] <= 8'h00;
memory0_reg[816 ] <= 8'h00;
memory0_reg[817 ] <= 8'h00;
memory0_reg[818 ] <= 8'h00;
memory0_reg[819 ] <= 8'h00;
memory0_reg[820 ] <= 8'h00;
memory0_reg[821 ] <= 8'h00;
memory0_reg[822 ] <= 8'h00;
memory0_reg[823 ] <= 8'h00;
memory0_reg[824 ] <= 8'h00;
memory0_reg[825 ] <= 8'h00;
memory0_reg[826 ] <= 8'h00;
memory0_reg[827 ] <= 8'h00;
memory0_reg[828 ] <= 8'h00;
memory0_reg[829 ] <= 8'h00;
memory0_reg[830 ] <= 8'h00;
memory0_reg[831 ] <= 8'h00;
memory0_reg[832 ] <= 8'h00;
memory0_reg[833 ] <= 8'h00;
memory0_reg[834 ] <= 8'h00;
memory0_reg[835 ] <= 8'h00;
memory0_reg[836 ] <= 8'h00;
memory0_reg[837 ] <= 8'h00;
memory0_reg[838 ] <= 8'h00;
memory0_reg[839 ] <= 8'h00;
memory0_reg[840 ] <= 8'h00;
memory0_reg[841 ] <= 8'h00;
memory0_reg[842 ] <= 8'h00;
memory0_reg[843 ] <= 8'h00;
memory0_reg[844 ] <= 8'h00;
memory0_reg[845 ] <= 8'h00;
memory0_reg[846 ] <= 8'h00;
memory0_reg[847 ] <= 8'h00;
memory0_reg[848 ] <= 8'h00;
memory0_reg[849 ] <= 8'h00;
memory0_reg[850 ] <= 8'h00;
memory0_reg[851 ] <= 8'h00;
memory0_reg[852 ] <= 8'h00;
memory0_reg[853 ] <= 8'h00;
memory0_reg[854 ] <= 8'h00;
memory0_reg[855 ] <= 8'h00;
memory0_reg[856 ] <= 8'h00;
memory0_reg[857 ] <= 8'h00;
memory0_reg[858 ] <= 8'h00;
memory0_reg[859 ] <= 8'h00;
memory0_reg[860 ] <= 8'h00;
memory0_reg[861 ] <= 8'h00;
memory0_reg[862 ] <= 8'h00;
memory0_reg[863 ] <= 8'h00;
memory0_reg[864 ] <= 8'h00;
memory0_reg[865 ] <= 8'h00;
memory0_reg[866 ] <= 8'h00;
memory0_reg[867 ] <= 8'h00;
memory0_reg[868 ] <= 8'h00;
memory0_reg[869 ] <= 8'h00;
memory0_reg[870 ] <= 8'h00;
memory0_reg[871 ] <= 8'h00;
memory0_reg[872 ] <= 8'h00;
memory0_reg[873 ] <= 8'h00;
memory0_reg[874 ] <= 8'h00;
memory0_reg[875 ] <= 8'h00;
memory0_reg[876 ] <= 8'h00;
memory0_reg[877 ] <= 8'h00;
memory0_reg[878 ] <= 8'h00;
memory0_reg[879 ] <= 8'h00;
memory0_reg[880 ] <= 8'h00;
memory0_reg[881 ] <= 8'h00;
memory0_reg[882 ] <= 8'h00;
memory0_reg[883 ] <= 8'h00;
memory0_reg[884 ] <= 8'h00;
memory0_reg[885 ] <= 8'h00;
memory0_reg[886 ] <= 8'h00;
memory0_reg[887 ] <= 8'h00;
memory0_reg[888 ] <= 8'h00;
memory0_reg[889 ] <= 8'h00;
memory0_reg[890 ] <= 8'h00;
memory0_reg[891 ] <= 8'h00;
memory0_reg[892 ] <= 8'h00;
memory0_reg[893 ] <= 8'h00;
memory0_reg[894 ] <= 8'h00;
memory0_reg[895 ] <= 8'h00;
memory0_reg[896 ] <= 8'h00;
memory0_reg[897 ] <= 8'h00;
memory0_reg[898 ] <= 8'h00;
memory0_reg[899 ] <= 8'h00;
memory0_reg[900 ] <= 8'h00;
memory0_reg[901 ] <= 8'h00;
memory0_reg[902 ] <= 8'h00;
memory0_reg[903 ] <= 8'h00;
memory0_reg[904 ] <= 8'h00;
memory0_reg[905 ] <= 8'h00;
memory0_reg[906 ] <= 8'h00;
memory0_reg[907 ] <= 8'h00;
memory0_reg[908 ] <= 8'h00;
memory0_reg[909 ] <= 8'h00;
memory0_reg[910 ] <= 8'h00;
memory0_reg[911 ] <= 8'h00;
memory0_reg[912 ] <= 8'h00;
memory0_reg[913 ] <= 8'h00;
memory0_reg[914 ] <= 8'h00;
memory0_reg[915 ] <= 8'h00;
memory0_reg[916 ] <= 8'h00;
memory0_reg[917 ] <= 8'h00;
memory0_reg[918 ] <= 8'h00;
memory0_reg[919 ] <= 8'h00;
memory0_reg[920 ] <= 8'h00;
memory0_reg[921 ] <= 8'h00;
memory0_reg[922 ] <= 8'h00;
memory0_reg[923 ] <= 8'h00;
memory0_reg[924 ] <= 8'h00;
memory0_reg[925 ] <= 8'h00;
memory0_reg[926 ] <= 8'h00;
memory0_reg[927 ] <= 8'h00;
memory0_reg[928 ] <= 8'h00;
memory0_reg[929 ] <= 8'h00;
memory0_reg[930 ] <= 8'h00;
memory0_reg[931 ] <= 8'h00;
memory0_reg[932 ] <= 8'h00;
memory0_reg[933 ] <= 8'h00;
memory0_reg[934 ] <= 8'h00;
memory0_reg[935 ] <= 8'h00;
memory0_reg[936 ] <= 8'h00;
memory0_reg[937 ] <= 8'h00;
memory0_reg[938 ] <= 8'h00;
memory0_reg[939 ] <= 8'h00;
memory0_reg[940 ] <= 8'h00;
memory0_reg[941 ] <= 8'h00;
memory0_reg[942 ] <= 8'h00;
memory0_reg[943 ] <= 8'h00;
memory0_reg[944 ] <= 8'h00;
memory0_reg[945 ] <= 8'h00;
memory0_reg[946 ] <= 8'h00;
memory0_reg[947 ] <= 8'h00;
memory0_reg[948 ] <= 8'h00;
memory0_reg[949 ] <= 8'h00;
memory0_reg[950 ] <= 8'h00;
memory0_reg[951 ] <= 8'h00;
memory0_reg[952 ] <= 8'h00;
memory0_reg[953 ] <= 8'h00;
memory0_reg[954 ] <= 8'h00;
memory0_reg[955 ] <= 8'h00;
memory0_reg[956 ] <= 8'h00;
memory0_reg[957 ] <= 8'h00;
memory0_reg[958 ] <= 8'h00;
memory0_reg[959 ] <= 8'h00;
memory0_reg[960 ] <= 8'h00;
memory0_reg[961 ] <= 8'h00;
memory0_reg[962 ] <= 8'h00;
memory0_reg[963 ] <= 8'h00;
memory0_reg[964 ] <= 8'h00;
memory0_reg[965 ] <= 8'h00;
memory0_reg[966 ] <= 8'h00;
memory0_reg[967 ] <= 8'h00;
memory0_reg[968 ] <= 8'h00;
memory0_reg[969 ] <= 8'h00;
memory0_reg[970 ] <= 8'h00;
memory0_reg[971 ] <= 8'h00;
memory0_reg[972 ] <= 8'h00;
memory0_reg[973 ] <= 8'h00;
memory0_reg[974 ] <= 8'h00;
memory0_reg[975 ] <= 8'h00;
memory0_reg[976 ] <= 8'h00;
memory0_reg[977 ] <= 8'h00;
memory0_reg[978 ] <= 8'h00;
memory0_reg[979 ] <= 8'h00;
memory0_reg[980 ] <= 8'h00;
memory0_reg[981 ] <= 8'h00;
memory0_reg[982 ] <= 8'h00;
memory0_reg[983 ] <= 8'h00;
memory0_reg[984 ] <= 8'h00;
memory0_reg[985 ] <= 8'h00;
memory0_reg[986 ] <= 8'h00;
memory0_reg[987 ] <= 8'h00;
memory0_reg[988 ] <= 8'h00;
memory0_reg[989 ] <= 8'h00;
memory0_reg[990 ] <= 8'h00;
memory0_reg[991 ] <= 8'h00;
memory0_reg[992 ] <= 8'h00;
memory0_reg[993 ] <= 8'h00;
memory0_reg[994 ] <= 8'h00;
memory0_reg[995 ] <= 8'h00;
memory0_reg[996 ] <= 8'h00;
memory0_reg[997 ] <= 8'h00;
memory0_reg[998 ] <= 8'h00;
memory0_reg[999 ] <= 8'h00;
memory0_reg[1000] <= 8'h00;
memory0_reg[1001] <= 8'h00;
memory0_reg[1002] <= 8'h00;
memory0_reg[1003] <= 8'h00;
memory0_reg[1004] <= 8'h00;
memory0_reg[1005] <= 8'h00;
memory0_reg[1006] <= 8'h00;
memory0_reg[1007] <= 8'h00;
memory0_reg[1008] <= 8'h00;
memory0_reg[1009] <= 8'h00;
memory0_reg[1010] <= 8'h00;
memory0_reg[1011] <= 8'h00;
memory0_reg[1012] <= 8'h00;
memory0_reg[1013] <= 8'h00;
memory0_reg[1014] <= 8'h00;
memory0_reg[1015] <= 8'h00;
memory0_reg[1016] <= 8'h00;
memory0_reg[1017] <= 8'h00;
memory0_reg[1018] <= 8'h00;
memory0_reg[1019] <= 8'h00;
memory0_reg[1020] <= 8'h00;
memory0_reg[1021] <= 8'h00;
memory0_reg[1022] <= 8'h00;
memory0_reg[1023] <= 8'h00;

// Memory 1

memory1_reg[0   ] <= 8'h00;
memory1_reg[1   ] <= 8'h00;
memory1_reg[2   ] <= 8'h00;
memory1_reg[3   ] <= 8'h00;
memory1_reg[4   ] <= 8'h00;
memory1_reg[5   ] <= 8'h00;
memory1_reg[6   ] <= 8'h00;
memory1_reg[7   ] <= 8'h00;
memory1_reg[8   ] <= 8'h00;
memory1_reg[9   ] <= 8'h00;
memory1_reg[10  ] <= 8'h02;
memory1_reg[11  ] <= 8'h00;
memory1_reg[12  ] <= 8'h00;
memory1_reg[13  ] <= 8'h00;
memory1_reg[14  ] <= 8'h00;
memory1_reg[15  ] <= 8'h00;
memory1_reg[16  ] <= 8'h00;
memory1_reg[17  ] <= 8'h0A;
memory1_reg[18  ] <= 8'h00;
memory1_reg[19  ] <= 8'h00;
memory1_reg[20  ] <= 8'h00;
memory1_reg[21  ] <= 8'h00;
memory1_reg[22  ] <= 8'h00;
memory1_reg[23  ] <= 8'h00;
memory1_reg[24  ] <= 8'h00;
memory1_reg[25  ] <= 8'h00;
memory1_reg[26  ] <= 8'h00;
memory1_reg[27  ] <= 8'h00;
memory1_reg[28  ] <= 8'h02;
memory1_reg[29  ] <= 8'h00;
memory1_reg[30  ] <= 8'h00;
memory1_reg[31  ] <= 8'h00;
memory1_reg[32  ] <= 8'h00;
memory1_reg[33  ] <= 8'h00;
memory1_reg[34  ] <= 8'h00;
memory1_reg[35  ] <= 8'h0A;
memory1_reg[36  ] <= 8'h00;
memory1_reg[37  ] <= 8'h00;
memory1_reg[38  ] <= 8'h00;
memory1_reg[39  ] <= 8'h00;
memory1_reg[40  ] <= 8'h00;
memory1_reg[41  ] <= 8'h00;
memory1_reg[42  ] <= 8'h00;
memory1_reg[43  ] <= 8'h00;
memory1_reg[44  ] <= 8'h00;
memory1_reg[45  ] <= 8'h00;
memory1_reg[46  ] <= 8'h02;
memory1_reg[47  ] <= 8'h00;
memory1_reg[48  ] <= 8'h00;
memory1_reg[49  ] <= 8'h00;
memory1_reg[50  ] <= 8'h00;
memory1_reg[51  ] <= 8'h00;
memory1_reg[52  ] <= 8'h00;
memory1_reg[53  ] <= 8'h06;
memory1_reg[54  ] <= 8'h00;
memory1_reg[55  ] <= 8'h00;
memory1_reg[56  ] <= 8'h00;
memory1_reg[57  ] <= 8'h00;
memory1_reg[58  ] <= 8'h00;
memory1_reg[59  ] <= 8'h00;
memory1_reg[60  ] <= 8'h00;
memory1_reg[61  ] <= 8'h00;
memory1_reg[62  ] <= 8'h00;
memory1_reg[63  ] <= 8'h00;
memory1_reg[64  ] <= 8'h00;
memory1_reg[65  ] <= 8'h00;
memory1_reg[66  ] <= 8'h02;
memory1_reg[67  ] <= 8'h00;
memory1_reg[68  ] <= 8'h00;
memory1_reg[69  ] <= 8'h00;
memory1_reg[70  ] <= 8'h00;
memory1_reg[71  ] <= 8'h00;
memory1_reg[72  ] <= 8'h00;
memory1_reg[73  ] <= 8'h0A;
memory1_reg[74  ] <= 8'h00;
memory1_reg[75  ] <= 8'h00;
memory1_reg[76  ] <= 8'h00;
memory1_reg[77  ] <= 8'h00;
memory1_reg[78  ] <= 8'h00;
memory1_reg[79  ] <= 8'h00;
memory1_reg[80  ] <= 8'h00;
memory1_reg[81  ] <= 8'h00;
memory1_reg[82  ] <= 8'h00;
memory1_reg[83  ] <= 8'h00;
memory1_reg[84  ] <= 8'h02;
memory1_reg[85  ] <= 8'h00;
memory1_reg[86  ] <= 8'h00;
memory1_reg[87  ] <= 8'h00;
memory1_reg[88  ] <= 8'h00;
memory1_reg[89  ] <= 8'h00;
memory1_reg[90  ] <= 8'h00;
memory1_reg[91  ] <= 8'h0A;
memory1_reg[92  ] <= 8'h00;
memory1_reg[93  ] <= 8'h00;
memory1_reg[94  ] <= 8'h00;
memory1_reg[95  ] <= 8'h00;
memory1_reg[96  ] <= 8'h00;
memory1_reg[97  ] <= 8'h00;
memory1_reg[98  ] <= 8'h00;
memory1_reg[99  ] <= 8'h00;
memory1_reg[100 ] <= 8'h00;
memory1_reg[101 ] <= 8'h00;
memory1_reg[102 ] <= 8'h02;
memory1_reg[103 ] <= 8'h00;
memory1_reg[104 ] <= 8'h00;
memory1_reg[105 ] <= 8'h00;
memory1_reg[106 ] <= 8'h00;
memory1_reg[107 ] <= 8'h00;
memory1_reg[108 ] <= 8'h00;
memory1_reg[109 ] <= 8'h06;
memory1_reg[110 ] <= 8'h00;
memory1_reg[111 ] <= 8'h00;
memory1_reg[112 ] <= 8'h00;
memory1_reg[113 ] <= 8'h00;
memory1_reg[114 ] <= 8'h00;
memory1_reg[115 ] <= 8'h00;
memory1_reg[116 ] <= 8'h00;
memory1_reg[117 ] <= 8'h00;
memory1_reg[118 ] <= 8'h00;
memory1_reg[119 ] <= 8'h00;
memory1_reg[120 ] <= 8'h00;
memory1_reg[121 ] <= 8'h00;
memory1_reg[122 ] <= 8'h02;
memory1_reg[123 ] <= 8'h00;
memory1_reg[124 ] <= 8'h00;
memory1_reg[125 ] <= 8'h00;
memory1_reg[126 ] <= 8'h00;
memory1_reg[127 ] <= 8'h00;
memory1_reg[128 ] <= 8'h00;
memory1_reg[129 ] <= 8'h0A;
memory1_reg[130 ] <= 8'h00;
memory1_reg[131 ] <= 8'h00;
memory1_reg[132 ] <= 8'h00;
memory1_reg[133 ] <= 8'h00;
memory1_reg[134 ] <= 8'h00;
memory1_reg[135 ] <= 8'h00;
memory1_reg[136 ] <= 8'h00;
memory1_reg[137 ] <= 8'h00;
memory1_reg[138 ] <= 8'h00;
memory1_reg[139 ] <= 8'h00;
memory1_reg[140 ] <= 8'h02;
memory1_reg[141 ] <= 8'h00;
memory1_reg[142 ] <= 8'h00;
memory1_reg[143 ] <= 8'h00;
memory1_reg[144 ] <= 8'h00;
memory1_reg[145 ] <= 8'h00;
memory1_reg[146 ] <= 8'h00;
memory1_reg[147 ] <= 8'h0A;
memory1_reg[148 ] <= 8'h00;
memory1_reg[149 ] <= 8'h00;
memory1_reg[150 ] <= 8'h00;
memory1_reg[151 ] <= 8'h00;
memory1_reg[152 ] <= 8'h00;
memory1_reg[153 ] <= 8'h00;
memory1_reg[154 ] <= 8'h00;
memory1_reg[155 ] <= 8'h00;
memory1_reg[156 ] <= 8'h00;
memory1_reg[157 ] <= 8'h00;
memory1_reg[158 ] <= 8'h02;
memory1_reg[159 ] <= 8'h00;
memory1_reg[160 ] <= 8'h00;
memory1_reg[161 ] <= 8'h00;
memory1_reg[162 ] <= 8'h00;
memory1_reg[163 ] <= 8'h00;
memory1_reg[164 ] <= 8'h00;
memory1_reg[165 ] <= 8'h06;
memory1_reg[166 ] <= 8'h00;
memory1_reg[167 ] <= 8'h00;
memory1_reg[168 ] <= 8'h00;
memory1_reg[169 ] <= 8'h00;
memory1_reg[170 ] <= 8'h00;
memory1_reg[171 ] <= 8'h00;
memory1_reg[172 ] <= 8'h00;
memory1_reg[173 ] <= 8'h00;
memory1_reg[174 ] <= 8'h00;
memory1_reg[175 ] <= 8'h00;
memory1_reg[176 ] <= 8'h00;
memory1_reg[177 ] <= 8'h02;
memory1_reg[178 ] <= 8'h00;
memory1_reg[179 ] <= 8'h00;
memory1_reg[180 ] <= 8'h00;
memory1_reg[181 ] <= 8'h00;
memory1_reg[182 ] <= 8'h00;
memory1_reg[183 ] <= 8'h00;
memory1_reg[184 ] <= 8'h00;
memory1_reg[185 ] <= 8'h00;
memory1_reg[186 ] <= 8'h00;
memory1_reg[187 ] <= 8'h02;
memory1_reg[188 ] <= 8'h00;
memory1_reg[189 ] <= 8'h00;
memory1_reg[190 ] <= 8'h00;
memory1_reg[191 ] <= 8'h00;
memory1_reg[192 ] <= 8'h00;
memory1_reg[193 ] <= 8'h00;
memory1_reg[194 ] <= 8'h00;
memory1_reg[195 ] <= 8'h00;
memory1_reg[196 ] <= 8'h00;
memory1_reg[197 ] <= 8'h0E;
memory1_reg[198 ] <= 8'h00;
memory1_reg[199 ] <= 8'h00;
memory1_reg[200 ] <= 8'h00;
memory1_reg[201 ] <= 8'h00;
memory1_reg[202 ] <= 8'h00;
memory1_reg[203 ] <= 8'h00;
memory1_reg[204 ] <= 8'h00;
memory1_reg[205 ] <= 8'h00;
memory1_reg[206 ] <= 8'h00;
memory1_reg[207 ] <= 8'h00;
memory1_reg[208 ] <= 8'h00;
memory1_reg[209 ] <= 8'h00;
memory1_reg[210 ] <= 8'h00;
memory1_reg[211 ] <= 8'h00;
memory1_reg[212 ] <= 8'h00;
memory1_reg[213 ] <= 8'h00;
memory1_reg[214 ] <= 8'h00;
memory1_reg[215 ] <= 8'h00;
memory1_reg[216 ] <= 8'h00;
memory1_reg[217 ] <= 8'h00;
memory1_reg[218 ] <= 8'h00;
memory1_reg[219 ] <= 8'h00;
memory1_reg[220 ] <= 8'h00;
memory1_reg[221 ] <= 8'h00;
memory1_reg[222 ] <= 8'h00;
memory1_reg[223 ] <= 8'h00;
memory1_reg[224 ] <= 8'h00;
memory1_reg[225 ] <= 8'h00;
memory1_reg[226 ] <= 8'h00;
memory1_reg[227 ] <= 8'h00;
memory1_reg[228 ] <= 8'h00;
memory1_reg[229 ] <= 8'h00;
memory1_reg[230 ] <= 8'h00;
memory1_reg[231 ] <= 8'h00;
memory1_reg[232 ] <= 8'h00;
memory1_reg[233 ] <= 8'h00;
memory1_reg[234 ] <= 8'h00;
memory1_reg[235 ] <= 8'h00;
memory1_reg[236 ] <= 8'h00;
memory1_reg[237 ] <= 8'h00;
memory1_reg[238 ] <= 8'h00;
memory1_reg[239 ] <= 8'h00;
memory1_reg[240 ] <= 8'h00;
memory1_reg[241 ] <= 8'h00;
memory1_reg[242 ] <= 8'h00;
memory1_reg[243 ] <= 8'h00;
memory1_reg[244 ] <= 8'h00;
memory1_reg[245 ] <= 8'h00;
memory1_reg[246 ] <= 8'h00;
memory1_reg[247 ] <= 8'h00;
memory1_reg[248 ] <= 8'h00;
memory1_reg[249 ] <= 8'h00;
memory1_reg[250 ] <= 8'h00;
memory1_reg[251 ] <= 8'h00;
memory1_reg[252 ] <= 8'h00;
memory1_reg[253 ] <= 8'h00;
memory1_reg[254 ] <= 8'h00;
memory1_reg[255 ] <= 8'h00;
memory1_reg[256 ] <= 8'h00;
memory1_reg[257 ] <= 8'h00;
memory1_reg[258 ] <= 8'h00;
memory1_reg[259 ] <= 8'h00;
memory1_reg[260 ] <= 8'h00;
memory1_reg[261 ] <= 8'h00;
memory1_reg[262 ] <= 8'h00;
memory1_reg[263 ] <= 8'h02;
memory1_reg[264 ] <= 8'h00;
memory1_reg[265 ] <= 8'h00;
memory1_reg[266 ] <= 8'h00;
memory1_reg[267 ] <= 8'h00;
memory1_reg[268 ] <= 8'h00;
memory1_reg[269 ] <= 8'h00;
memory1_reg[270 ] <= 8'h02;
memory1_reg[271 ] <= 8'h00;
memory1_reg[272 ] <= 8'h00;
memory1_reg[273 ] <= 8'h00;
memory1_reg[274 ] <= 8'h00;
memory1_reg[275 ] <= 8'h00;
memory1_reg[276 ] <= 8'h00;
memory1_reg[277 ] <= 8'h02;
memory1_reg[278 ] <= 8'h00;
memory1_reg[279 ] <= 8'h00;
memory1_reg[280 ] <= 8'h00;
memory1_reg[281 ] <= 8'h00;
memory1_reg[282 ] <= 8'h00;
memory1_reg[283 ] <= 8'h00;
memory1_reg[284 ] <= 8'h02;
memory1_reg[285 ] <= 8'h00;
memory1_reg[286 ] <= 8'h00;
memory1_reg[287 ] <= 8'h00;
memory1_reg[288 ] <= 8'h00;
memory1_reg[289 ] <= 8'h00;
memory1_reg[290 ] <= 8'h00;
memory1_reg[291 ] <= 8'h02;
memory1_reg[292 ] <= 8'h00;
memory1_reg[293 ] <= 8'h00;
memory1_reg[294 ] <= 8'h00;
memory1_reg[295 ] <= 8'h00;
memory1_reg[296 ] <= 8'h00;
memory1_reg[297 ] <= 8'h00;
memory1_reg[298 ] <= 8'h02;
memory1_reg[299 ] <= 8'h00;
memory1_reg[300 ] <= 8'h00;
memory1_reg[301 ] <= 8'h00;
memory1_reg[302 ] <= 8'h00;
memory1_reg[303 ] <= 8'h00;
memory1_reg[304 ] <= 8'h00;
memory1_reg[305 ] <= 8'h02;
memory1_reg[306 ] <= 8'h00;
memory1_reg[307 ] <= 8'h00;
memory1_reg[308 ] <= 8'h00;
memory1_reg[309 ] <= 8'h00;
memory1_reg[310 ] <= 8'h00;
memory1_reg[311 ] <= 8'h00;
memory1_reg[312 ] <= 8'h02;
memory1_reg[313 ] <= 8'h00;
memory1_reg[314 ] <= 8'h00;
memory1_reg[315 ] <= 8'h00;
memory1_reg[316 ] <= 8'h00;
memory1_reg[317 ] <= 8'h00;
memory1_reg[318 ] <= 8'h00;
memory1_reg[319 ] <= 8'h06;
memory1_reg[320 ] <= 8'h00;
memory1_reg[321 ] <= 8'h01;
memory1_reg[322 ] <= 8'h00;
memory1_reg[323 ] <= 8'h00;
memory1_reg[324 ] <= 8'h00;
memory1_reg[325 ] <= 8'h00;
memory1_reg[326 ] <= 8'h00;
memory1_reg[327 ] <= 8'h00;
memory1_reg[328 ] <= 8'h02;
memory1_reg[329 ] <= 8'h01;
memory1_reg[330 ] <= 8'h00;
memory1_reg[331 ] <= 8'h00;
memory1_reg[332 ] <= 8'h00;
memory1_reg[333 ] <= 8'h00;
memory1_reg[334 ] <= 8'h00;
memory1_reg[335 ] <= 8'h00;
memory1_reg[336 ] <= 8'h02;
memory1_reg[337 ] <= 8'h01;
memory1_reg[338 ] <= 8'h00;
memory1_reg[339 ] <= 8'h00;
memory1_reg[340 ] <= 8'h00;
memory1_reg[341 ] <= 8'h00;
memory1_reg[342 ] <= 8'h00;
memory1_reg[343 ] <= 8'h00;
memory1_reg[344 ] <= 8'h02;
memory1_reg[345 ] <= 8'h00;
memory1_reg[346 ] <= 8'h00;
memory1_reg[347 ] <= 8'h0E;
memory1_reg[348 ] <= 8'h04;
memory1_reg[349 ] <= 8'h00;
memory1_reg[350 ] <= 8'h00;
memory1_reg[351 ] <= 8'h00;
memory1_reg[352 ] <= 8'h04;
memory1_reg[353 ] <= 8'h00;
memory1_reg[354 ] <= 8'h00;
memory1_reg[355 ] <= 8'h00;
memory1_reg[356 ] <= 8'h04;
memory1_reg[357 ] <= 8'h00;
memory1_reg[358 ] <= 8'h00;
memory1_reg[359 ] <= 8'h00;
memory1_reg[360 ] <= 8'h04;
memory1_reg[361 ] <= 8'h00;
memory1_reg[362 ] <= 8'h00;
memory1_reg[363 ] <= 8'h00;
memory1_reg[364 ] <= 8'h0C;
memory1_reg[365 ] <= 8'h00;
memory1_reg[366 ] <= 8'h00;
memory1_reg[367 ] <= 8'h00;
memory1_reg[368 ] <= 8'h01;
memory1_reg[369 ] <= 8'h06;
memory1_reg[370 ] <= 8'h00;
memory1_reg[371 ] <= 8'h00;
memory1_reg[372 ] <= 8'h00;
memory1_reg[373 ] <= 8'h00;
memory1_reg[374 ] <= 8'h00;
memory1_reg[375 ] <= 8'h06;
memory1_reg[376 ] <= 8'h00;
memory1_reg[377 ] <= 8'h00;
memory1_reg[378 ] <= 8'h00;
memory1_reg[379 ] <= 8'h06;
memory1_reg[380 ] <= 8'h00;
memory1_reg[381 ] <= 8'h00;
memory1_reg[382 ] <= 8'h00;
memory1_reg[383 ] <= 8'h06;
memory1_reg[384 ] <= 8'h00;
memory1_reg[385 ] <= 8'h01;
memory1_reg[386 ] <= 8'h00;
memory1_reg[387 ] <= 8'h00;
memory1_reg[388 ] <= 8'h00;
memory1_reg[389 ] <= 8'h00;
memory1_reg[390 ] <= 8'h00;
memory1_reg[391 ] <= 8'h00;
memory1_reg[392 ] <= 8'h02;
memory1_reg[393 ] <= 8'h01;
memory1_reg[394 ] <= 8'h00;
memory1_reg[395 ] <= 8'h00;
memory1_reg[396 ] <= 8'h00;
memory1_reg[397 ] <= 8'h00;
memory1_reg[398 ] <= 8'h00;
memory1_reg[399 ] <= 8'h00;
memory1_reg[400 ] <= 8'h02;
memory1_reg[401 ] <= 8'h01;
memory1_reg[402 ] <= 8'h00;
memory1_reg[403 ] <= 8'h00;
memory1_reg[404 ] <= 8'h00;
memory1_reg[405 ] <= 8'h00;
memory1_reg[406 ] <= 8'h00;
memory1_reg[407 ] <= 8'h00;
memory1_reg[408 ] <= 8'h0E;
memory1_reg[409 ] <= 8'h00;
memory1_reg[410 ] <= 8'h00;
memory1_reg[411 ] <= 8'h00;
memory1_reg[412 ] <= 8'h00;
memory1_reg[413 ] <= 8'h00;
memory1_reg[414 ] <= 8'h00;
memory1_reg[415 ] <= 8'h02;
memory1_reg[416 ] <= 8'h00;
memory1_reg[417 ] <= 8'h00;
memory1_reg[418 ] <= 8'h00;
memory1_reg[419 ] <= 8'h02;
memory1_reg[420 ] <= 8'h00;
memory1_reg[421 ] <= 8'h00;
memory1_reg[422 ] <= 8'h00;
memory1_reg[423 ] <= 8'h02;
memory1_reg[424 ] <= 8'h00;
memory1_reg[425 ] <= 8'h00;
memory1_reg[426 ] <= 8'h00;
memory1_reg[427 ] <= 8'h02;
memory1_reg[428 ] <= 8'h00;
memory1_reg[429 ] <= 8'h00;
memory1_reg[430 ] <= 8'h00;
memory1_reg[431 ] <= 8'h02;
memory1_reg[432 ] <= 8'h00;
memory1_reg[433 ] <= 8'h00;
memory1_reg[434 ] <= 8'h00;
memory1_reg[435 ] <= 8'h02;
memory1_reg[436 ] <= 8'h00;
memory1_reg[437 ] <= 8'h00;
memory1_reg[438 ] <= 8'h00;
memory1_reg[439 ] <= 8'h00;
memory1_reg[440 ] <= 8'h00;
memory1_reg[441 ] <= 8'h00;
memory1_reg[442 ] <= 8'h00;
memory1_reg[443 ] <= 8'h02;
memory1_reg[444 ] <= 8'h00;
memory1_reg[445 ] <= 8'h00;
memory1_reg[446 ] <= 8'h00;
memory1_reg[447 ] <= 8'h00;
memory1_reg[448 ] <= 8'h00;
memory1_reg[449 ] <= 8'h00;
memory1_reg[450 ] <= 8'h02;
memory1_reg[451 ] <= 8'h00;
memory1_reg[452 ] <= 8'h00;
memory1_reg[453 ] <= 8'h00;
memory1_reg[454 ] <= 8'h00;
memory1_reg[455 ] <= 8'h00;
memory1_reg[456 ] <= 8'h00;
memory1_reg[457 ] <= 8'h0A;
memory1_reg[458 ] <= 8'h00;
memory1_reg[459 ] <= 8'h00;
memory1_reg[460 ] <= 8'h02;
memory1_reg[461 ] <= 8'h00;
memory1_reg[462 ] <= 8'h00;
memory1_reg[463 ] <= 8'h02;
memory1_reg[464 ] <= 8'h00;
memory1_reg[465 ] <= 8'h00;
memory1_reg[466 ] <= 8'h02;
memory1_reg[467 ] <= 8'h00;
memory1_reg[468 ] <= 8'h00;
memory1_reg[469 ] <= 8'h02;
memory1_reg[470 ] <= 8'h00;
memory1_reg[471 ] <= 8'h00;
memory1_reg[472 ] <= 8'h06;
memory1_reg[473 ] <= 8'h00;
memory1_reg[474 ] <= 8'h00;
memory1_reg[475 ] <= 8'h00;
memory1_reg[476 ] <= 8'h01;
memory1_reg[477 ] <= 8'h02;
memory1_reg[478 ] <= 8'h01;
memory1_reg[479 ] <= 8'h02;
memory1_reg[480 ] <= 8'h01;
memory1_reg[481 ] <= 8'h0A;
memory1_reg[482 ] <= 8'h01;
memory1_reg[483 ] <= 8'h02;
memory1_reg[484 ] <= 8'h01;
memory1_reg[485 ] <= 8'h02;
memory1_reg[486 ] <= 8'h01;
memory1_reg[487 ] <= 8'h0A;
memory1_reg[488 ] <= 8'h01;
memory1_reg[489 ] <= 8'h02;
memory1_reg[490 ] <= 8'h01;
memory1_reg[491 ] <= 8'h02;
memory1_reg[492 ] <= 8'h01;
memory1_reg[493 ] <= 8'h0A;
memory1_reg[494 ] <= 8'h01;
memory1_reg[495 ] <= 8'h02;
memory1_reg[496 ] <= 8'h01;
memory1_reg[497 ] <= 8'h02;
memory1_reg[498 ] <= 8'h01;
memory1_reg[499 ] <= 8'h06;
memory1_reg[500 ] <= 8'h00;
memory1_reg[501 ] <= 8'h00;
memory1_reg[502 ] <= 8'h00;
memory1_reg[503 ] <= 8'h00;
memory1_reg[504 ] <= 8'h00;
memory1_reg[505 ] <= 8'h00;
memory1_reg[506 ] <= 8'h00;
memory1_reg[507 ] <= 8'h00;
memory1_reg[508 ] <= 8'h00;
memory1_reg[509 ] <= 8'h00;
memory1_reg[510 ] <= 8'h00;
memory1_reg[511 ] <= 8'h00;
memory1_reg[512 ] <= 8'h01;
memory1_reg[513 ] <= 8'h02;
memory1_reg[514 ] <= 8'h01;
memory1_reg[515 ] <= 8'h02;
memory1_reg[516 ] <= 8'h01;
memory1_reg[517 ] <= 8'h0A;
memory1_reg[518 ] <= 8'h01;
memory1_reg[519 ] <= 8'h02;
memory1_reg[520 ] <= 8'h01;
memory1_reg[521 ] <= 8'h02;
memory1_reg[522 ] <= 8'h01;
memory1_reg[523 ] <= 8'h0A;
memory1_reg[524 ] <= 8'h01;
memory1_reg[525 ] <= 8'h02;
memory1_reg[526 ] <= 8'h01;
memory1_reg[527 ] <= 8'h02;
memory1_reg[528 ] <= 8'h01;
memory1_reg[529 ] <= 8'h0A;
memory1_reg[530 ] <= 8'h01;
memory1_reg[531 ] <= 8'h02;
memory1_reg[532 ] <= 8'h01;
memory1_reg[533 ] <= 8'h02;
memory1_reg[534 ] <= 8'h01;
memory1_reg[535 ] <= 8'h06;
memory1_reg[536 ] <= 8'h00;
memory1_reg[537 ] <= 8'h00;
memory1_reg[538 ] <= 8'h00;
memory1_reg[539 ] <= 8'h02;
memory1_reg[540 ] <= 8'h00;
memory1_reg[541 ] <= 8'h00;
memory1_reg[542 ] <= 8'h06;
memory1_reg[543 ] <= 8'h00;
memory1_reg[544 ] <= 8'h00;
memory1_reg[545 ] <= 8'h00;
memory1_reg[546 ] <= 8'h00;
memory1_reg[547 ] <= 8'h00;
memory1_reg[548 ] <= 8'h00;
memory1_reg[549 ] <= 8'h06;
memory1_reg[550 ] <= 8'h00;
memory1_reg[551 ] <= 8'h00;
memory1_reg[552 ] <= 8'h00;
memory1_reg[553 ] <= 8'h00;
memory1_reg[554 ] <= 8'h02;
memory1_reg[555 ] <= 8'h00;
memory1_reg[556 ] <= 8'h00;
memory1_reg[557 ] <= 8'h02;
memory1_reg[558 ] <= 8'h00;
memory1_reg[559 ] <= 8'h00;
memory1_reg[560 ] <= 8'h02;
memory1_reg[561 ] <= 8'h00;
memory1_reg[562 ] <= 8'h00;
memory1_reg[563 ] <= 8'h00;
memory1_reg[564 ] <= 8'h00;
memory1_reg[565 ] <= 8'h00;
memory1_reg[566 ] <= 8'h00;
memory1_reg[567 ] <= 8'h00;
memory1_reg[568 ] <= 8'h00;
memory1_reg[569 ] <= 8'h02;
memory1_reg[570 ] <= 8'h00;
memory1_reg[571 ] <= 8'h00;
memory1_reg[572 ] <= 8'h00;
memory1_reg[573 ] <= 8'h00;
memory1_reg[574 ] <= 8'h00;
memory1_reg[575 ] <= 8'h00;
memory1_reg[576 ] <= 8'h00;
memory1_reg[577 ] <= 8'h00;
memory1_reg[578 ] <= 8'h02;
memory1_reg[579 ] <= 8'h00;
memory1_reg[580 ] <= 8'h00;
memory1_reg[581 ] <= 8'h00;
memory1_reg[582 ] <= 8'h00;
memory1_reg[583 ] <= 8'h00;
memory1_reg[584 ] <= 8'h00;
memory1_reg[585 ] <= 8'h00;
memory1_reg[586 ] <= 8'h02;
memory1_reg[587 ] <= 8'h00;
memory1_reg[588 ] <= 8'h00;
memory1_reg[589 ] <= 8'h00;
memory1_reg[590 ] <= 8'h00;
memory1_reg[591 ] <= 8'h00;
memory1_reg[592 ] <= 8'h00;
memory1_reg[593 ] <= 8'h00;
memory1_reg[594 ] <= 8'h00;
memory1_reg[595 ] <= 8'h06;
memory1_reg[596 ] <= 8'h00;
memory1_reg[597 ] <= 8'h00;
memory1_reg[598 ] <= 8'h00;
memory1_reg[599 ] <= 8'h02;
memory1_reg[600 ] <= 8'h00;
memory1_reg[601 ] <= 8'h00;
memory1_reg[602 ] <= 8'h00;
memory1_reg[603 ] <= 8'h00;
memory1_reg[604 ] <= 8'h00;
memory1_reg[605 ] <= 8'h00;
memory1_reg[606 ] <= 8'h00;
memory1_reg[607 ] <= 8'h02;
memory1_reg[608 ] <= 8'h00;
memory1_reg[609 ] <= 8'h00;
memory1_reg[610 ] <= 8'h00;
memory1_reg[611 ] <= 8'h00;
memory1_reg[612 ] <= 8'h00;
memory1_reg[613 ] <= 8'h00;
memory1_reg[614 ] <= 8'h02;
memory1_reg[615 ] <= 8'h00;
memory1_reg[616 ] <= 8'h00;
memory1_reg[617 ] <= 8'h00;
memory1_reg[618 ] <= 8'h00;
memory1_reg[619 ] <= 8'h00;
memory1_reg[620 ] <= 8'h00;
memory1_reg[621 ] <= 8'h02;
memory1_reg[622 ] <= 8'h01;
memory1_reg[623 ] <= 8'h00;
memory1_reg[624 ] <= 8'h00;
memory1_reg[625 ] <= 8'h00;
memory1_reg[626 ] <= 8'h00;
memory1_reg[627 ] <= 8'h00;
memory1_reg[628 ] <= 8'h00;
memory1_reg[629 ] <= 8'h06;
memory1_reg[630 ] <= 8'h00;
memory1_reg[631 ] <= 8'h00;
memory1_reg[632 ] <= 8'h00;
memory1_reg[633 ] <= 8'h00;
memory1_reg[634 ] <= 8'h00;
memory1_reg[635 ] <= 8'h02;
memory1_reg[636 ] <= 8'h00;
memory1_reg[637 ] <= 8'h00;
memory1_reg[638 ] <= 8'h00;
memory1_reg[639 ] <= 8'h00;
memory1_reg[640 ] <= 8'h02;
memory1_reg[641 ] <= 8'h00;
memory1_reg[642 ] <= 8'h00;
memory1_reg[643 ] <= 8'h00;
memory1_reg[644 ] <= 8'h00;
memory1_reg[645 ] <= 8'h02;
memory1_reg[646 ] <= 8'h01;
memory1_reg[647 ] <= 8'h00;
memory1_reg[648 ] <= 8'h00;
memory1_reg[649 ] <= 8'h00;
memory1_reg[650 ] <= 8'h00;
memory1_reg[651 ] <= 8'h06;
memory1_reg[652 ] <= 8'h00;
memory1_reg[653 ] <= 8'h00;
memory1_reg[654 ] <= 8'h00;
memory1_reg[655 ] <= 8'h02;
memory1_reg[656 ] <= 8'h00;
memory1_reg[657 ] <= 8'h00;
memory1_reg[658 ] <= 8'h00;
memory1_reg[659 ] <= 8'h00;
memory1_reg[660 ] <= 8'h00;
memory1_reg[661 ] <= 8'h00;
memory1_reg[662 ] <= 8'h00;
memory1_reg[663 ] <= 8'h02;
memory1_reg[664 ] <= 8'h00;
memory1_reg[665 ] <= 8'h00;
memory1_reg[666 ] <= 8'h00;
memory1_reg[667 ] <= 8'h00;
memory1_reg[668 ] <= 8'h00;
memory1_reg[669 ] <= 8'h00;
memory1_reg[670 ] <= 8'h00;
memory1_reg[671 ] <= 8'h02;
memory1_reg[672 ] <= 8'h00;
memory1_reg[673 ] <= 8'h00;
memory1_reg[674 ] <= 8'h00;
memory1_reg[675 ] <= 8'h00;
memory1_reg[676 ] <= 8'h00;
memory1_reg[677 ] <= 8'h00;
memory1_reg[678 ] <= 8'h02;
memory1_reg[679 ] <= 8'h01;
memory1_reg[680 ] <= 8'h00;
memory1_reg[681 ] <= 8'h00;
memory1_reg[682 ] <= 8'h00;
memory1_reg[683 ] <= 8'h00;
memory1_reg[684 ] <= 8'h00;
memory1_reg[685 ] <= 8'h00;
memory1_reg[686 ] <= 8'h06;
memory1_reg[687 ] <= 8'h00;
memory1_reg[688 ] <= 8'h00;
memory1_reg[689 ] <= 8'h00;
memory1_reg[690 ] <= 8'h00;
memory1_reg[691 ] <= 8'h00;
memory1_reg[692 ] <= 8'h00;
memory1_reg[693 ] <= 8'h00;
memory1_reg[694 ] <= 8'h00;
memory1_reg[695 ] <= 8'h06;
memory1_reg[696 ] <= 8'h00;
memory1_reg[697 ] <= 8'h00;
memory1_reg[698 ] <= 8'h00;
memory1_reg[699 ] <= 8'h02;
memory1_reg[700 ] <= 8'h00;
memory1_reg[701 ] <= 8'h00;
memory1_reg[702 ] <= 8'h00;
memory1_reg[703 ] <= 8'h0A;
memory1_reg[704 ] <= 8'h00;
memory1_reg[705 ] <= 8'h00;
memory1_reg[706 ] <= 8'h00;
memory1_reg[707 ] <= 8'h0E;
memory1_reg[708 ] <= 8'h00;
memory1_reg[709 ] <= 8'h00;
memory1_reg[710 ] <= 8'h00;
memory1_reg[711 ] <= 8'h00;
memory1_reg[712 ] <= 8'h00;
memory1_reg[713 ] <= 8'h00;
memory1_reg[714 ] <= 8'h00;
memory1_reg[715 ] <= 8'h00;
memory1_reg[716 ] <= 8'h00;
memory1_reg[717 ] <= 8'h00;
memory1_reg[718 ] <= 8'h00;
memory1_reg[719 ] <= 8'h00;
memory1_reg[720 ] <= 8'h00;
memory1_reg[721 ] <= 8'h00;
memory1_reg[722 ] <= 8'h00;
memory1_reg[723 ] <= 8'h00;
memory1_reg[724 ] <= 8'h00;
memory1_reg[725 ] <= 8'h00;
memory1_reg[726 ] <= 8'h00;
memory1_reg[727 ] <= 8'h00;
memory1_reg[728 ] <= 8'h00;
memory1_reg[729 ] <= 8'h00;
memory1_reg[730 ] <= 8'h00;
memory1_reg[731 ] <= 8'h00;
memory1_reg[732 ] <= 8'h00;
memory1_reg[733 ] <= 8'h00;
memory1_reg[734 ] <= 8'h00;
memory1_reg[735 ] <= 8'h00;
memory1_reg[736 ] <= 8'h00;
memory1_reg[737 ] <= 8'h00;
memory1_reg[738 ] <= 8'h00;
memory1_reg[739 ] <= 8'h00;
memory1_reg[740 ] <= 8'h00;
memory1_reg[741 ] <= 8'h00;
memory1_reg[742 ] <= 8'h00;
memory1_reg[743 ] <= 8'h00;
memory1_reg[744 ] <= 8'h00;
memory1_reg[745 ] <= 8'h00;
memory1_reg[746 ] <= 8'h00;
memory1_reg[747 ] <= 8'h00;
memory1_reg[748 ] <= 8'h00;
memory1_reg[749 ] <= 8'h00;
memory1_reg[750 ] <= 8'h00;
memory1_reg[751 ] <= 8'h00;
memory1_reg[752 ] <= 8'h00;
memory1_reg[753 ] <= 8'h00;
memory1_reg[754 ] <= 8'h00;
memory1_reg[755 ] <= 8'h00;
memory1_reg[756 ] <= 8'h00;
memory1_reg[757 ] <= 8'h00;
memory1_reg[758 ] <= 8'h00;
memory1_reg[759 ] <= 8'h00;
memory1_reg[760 ] <= 8'h00;
memory1_reg[761 ] <= 8'h00;
memory1_reg[762 ] <= 8'h00;
memory1_reg[763 ] <= 8'h00;
memory1_reg[764 ] <= 8'h00;
memory1_reg[765 ] <= 8'h00;
memory1_reg[766 ] <= 8'h00;
memory1_reg[767 ] <= 8'h00;
memory1_reg[768 ] <= 8'h00;
memory1_reg[769 ] <= 8'h00;
memory1_reg[770 ] <= 8'h00;
memory1_reg[771 ] <= 8'h00;
memory1_reg[772 ] <= 8'h00;
memory1_reg[773 ] <= 8'h00;
memory1_reg[774 ] <= 8'h00;
memory1_reg[775 ] <= 8'h00;
memory1_reg[776 ] <= 8'h00;
memory1_reg[777 ] <= 8'h00;
memory1_reg[778 ] <= 8'h00;
memory1_reg[779 ] <= 8'h00;
memory1_reg[780 ] <= 8'h00;
memory1_reg[781 ] <= 8'h00;
memory1_reg[782 ] <= 8'h00;
memory1_reg[783 ] <= 8'h00;
memory1_reg[784 ] <= 8'h00;
memory1_reg[785 ] <= 8'h00;
memory1_reg[786 ] <= 8'h00;
memory1_reg[787 ] <= 8'h00;
memory1_reg[788 ] <= 8'h00;
memory1_reg[789 ] <= 8'h00;
memory1_reg[790 ] <= 8'h00;
memory1_reg[791 ] <= 8'h00;
memory1_reg[792 ] <= 8'h00;
memory1_reg[793 ] <= 8'h00;
memory1_reg[794 ] <= 8'h00;
memory1_reg[795 ] <= 8'h00;
memory1_reg[796 ] <= 8'h00;
memory1_reg[797 ] <= 8'h00;
memory1_reg[798 ] <= 8'h00;
memory1_reg[799 ] <= 8'h00;
memory1_reg[800 ] <= 8'h00;
memory1_reg[801 ] <= 8'h00;
memory1_reg[802 ] <= 8'h00;
memory1_reg[803 ] <= 8'h00;
memory1_reg[804 ] <= 8'h00;
memory1_reg[805 ] <= 8'h00;
memory1_reg[806 ] <= 8'h00;
memory1_reg[807 ] <= 8'h00;
memory1_reg[808 ] <= 8'h00;
memory1_reg[809 ] <= 8'h00;
memory1_reg[810 ] <= 8'h00;
memory1_reg[811 ] <= 8'h00;
memory1_reg[812 ] <= 8'h00;
memory1_reg[813 ] <= 8'h00;
memory1_reg[814 ] <= 8'h00;
memory1_reg[815 ] <= 8'h00;
memory1_reg[816 ] <= 8'h00;
memory1_reg[817 ] <= 8'h00;
memory1_reg[818 ] <= 8'h00;
memory1_reg[819 ] <= 8'h00;
memory1_reg[820 ] <= 8'h00;
memory1_reg[821 ] <= 8'h00;
memory1_reg[822 ] <= 8'h00;
memory1_reg[823 ] <= 8'h00;
memory1_reg[824 ] <= 8'h00;
memory1_reg[825 ] <= 8'h00;
memory1_reg[826 ] <= 8'h00;
memory1_reg[827 ] <= 8'h00;
memory1_reg[828 ] <= 8'h00;
memory1_reg[829 ] <= 8'h00;
memory1_reg[830 ] <= 8'h00;
memory1_reg[831 ] <= 8'h00;
memory1_reg[832 ] <= 8'h00;
memory1_reg[833 ] <= 8'h00;
memory1_reg[834 ] <= 8'h00;
memory1_reg[835 ] <= 8'h00;
memory1_reg[836 ] <= 8'h00;
memory1_reg[837 ] <= 8'h00;
memory1_reg[838 ] <= 8'h00;
memory1_reg[839 ] <= 8'h00;
memory1_reg[840 ] <= 8'h00;
memory1_reg[841 ] <= 8'h00;
memory1_reg[842 ] <= 8'h00;
memory1_reg[843 ] <= 8'h00;
memory1_reg[844 ] <= 8'h00;
memory1_reg[845 ] <= 8'h00;
memory1_reg[846 ] <= 8'h00;
memory1_reg[847 ] <= 8'h00;
memory1_reg[848 ] <= 8'h00;
memory1_reg[849 ] <= 8'h00;
memory1_reg[850 ] <= 8'h00;
memory1_reg[851 ] <= 8'h00;
memory1_reg[852 ] <= 8'h00;
memory1_reg[853 ] <= 8'h00;
memory1_reg[854 ] <= 8'h00;
memory1_reg[855 ] <= 8'h00;
memory1_reg[856 ] <= 8'h00;
memory1_reg[857 ] <= 8'h00;
memory1_reg[858 ] <= 8'h00;
memory1_reg[859 ] <= 8'h00;
memory1_reg[860 ] <= 8'h00;
memory1_reg[861 ] <= 8'h00;
memory1_reg[862 ] <= 8'h00;
memory1_reg[863 ] <= 8'h00;
memory1_reg[864 ] <= 8'h00;
memory1_reg[865 ] <= 8'h00;
memory1_reg[866 ] <= 8'h00;
memory1_reg[867 ] <= 8'h00;
memory1_reg[868 ] <= 8'h00;
memory1_reg[869 ] <= 8'h00;
memory1_reg[870 ] <= 8'h00;
memory1_reg[871 ] <= 8'h00;
memory1_reg[872 ] <= 8'h00;
memory1_reg[873 ] <= 8'h00;
memory1_reg[874 ] <= 8'h00;
memory1_reg[875 ] <= 8'h00;
memory1_reg[876 ] <= 8'h00;
memory1_reg[877 ] <= 8'h00;
memory1_reg[878 ] <= 8'h00;
memory1_reg[879 ] <= 8'h00;
memory1_reg[880 ] <= 8'h00;
memory1_reg[881 ] <= 8'h00;
memory1_reg[882 ] <= 8'h00;
memory1_reg[883 ] <= 8'h00;
memory1_reg[884 ] <= 8'h00;
memory1_reg[885 ] <= 8'h00;
memory1_reg[886 ] <= 8'h00;
memory1_reg[887 ] <= 8'h00;
memory1_reg[888 ] <= 8'h00;
memory1_reg[889 ] <= 8'h00;
memory1_reg[890 ] <= 8'h00;
memory1_reg[891 ] <= 8'h00;
memory1_reg[892 ] <= 8'h00;
memory1_reg[893 ] <= 8'h00;
memory1_reg[894 ] <= 8'h00;
memory1_reg[895 ] <= 8'h00;
memory1_reg[896 ] <= 8'h00;
memory1_reg[897 ] <= 8'h00;
memory1_reg[898 ] <= 8'h00;
memory1_reg[899 ] <= 8'h00;
memory1_reg[900 ] <= 8'h00;
memory1_reg[901 ] <= 8'h00;
memory1_reg[902 ] <= 8'h00;
memory1_reg[903 ] <= 8'h00;
memory1_reg[904 ] <= 8'h00;
memory1_reg[905 ] <= 8'h00;
memory1_reg[906 ] <= 8'h00;
memory1_reg[907 ] <= 8'h00;
memory1_reg[908 ] <= 8'h00;
memory1_reg[909 ] <= 8'h00;
memory1_reg[910 ] <= 8'h00;
memory1_reg[911 ] <= 8'h00;
memory1_reg[912 ] <= 8'h00;
memory1_reg[913 ] <= 8'h00;
memory1_reg[914 ] <= 8'h00;
memory1_reg[915 ] <= 8'h00;
memory1_reg[916 ] <= 8'h00;
memory1_reg[917 ] <= 8'h00;
memory1_reg[918 ] <= 8'h00;
memory1_reg[919 ] <= 8'h00;
memory1_reg[920 ] <= 8'h00;
memory1_reg[921 ] <= 8'h00;
memory1_reg[922 ] <= 8'h00;
memory1_reg[923 ] <= 8'h00;
memory1_reg[924 ] <= 8'h00;
memory1_reg[925 ] <= 8'h00;
memory1_reg[926 ] <= 8'h00;
memory1_reg[927 ] <= 8'h00;
memory1_reg[928 ] <= 8'h00;
memory1_reg[929 ] <= 8'h00;
memory1_reg[930 ] <= 8'h00;
memory1_reg[931 ] <= 8'h00;
memory1_reg[932 ] <= 8'h00;
memory1_reg[933 ] <= 8'h00;
memory1_reg[934 ] <= 8'h00;
memory1_reg[935 ] <= 8'h00;
memory1_reg[936 ] <= 8'h00;
memory1_reg[937 ] <= 8'h00;
memory1_reg[938 ] <= 8'h00;
memory1_reg[939 ] <= 8'h00;
memory1_reg[940 ] <= 8'h00;
memory1_reg[941 ] <= 8'h00;
memory1_reg[942 ] <= 8'h00;
memory1_reg[943 ] <= 8'h00;
memory1_reg[944 ] <= 8'h00;
memory1_reg[945 ] <= 8'h00;
memory1_reg[946 ] <= 8'h00;
memory1_reg[947 ] <= 8'h00;
memory1_reg[948 ] <= 8'h00;
memory1_reg[949 ] <= 8'h00;
memory1_reg[950 ] <= 8'h00;
memory1_reg[951 ] <= 8'h00;
memory1_reg[952 ] <= 8'h00;
memory1_reg[953 ] <= 8'h00;
memory1_reg[954 ] <= 8'h00;
memory1_reg[955 ] <= 8'h00;
memory1_reg[956 ] <= 8'h00;
memory1_reg[957 ] <= 8'h00;
memory1_reg[958 ] <= 8'h00;
memory1_reg[959 ] <= 8'h00;
memory1_reg[960 ] <= 8'h00;
memory1_reg[961 ] <= 8'h00;
memory1_reg[962 ] <= 8'h00;
memory1_reg[963 ] <= 8'h00;
memory1_reg[964 ] <= 8'h00;
memory1_reg[965 ] <= 8'h00;
memory1_reg[966 ] <= 8'h00;
memory1_reg[967 ] <= 8'h00;
memory1_reg[968 ] <= 8'h00;
memory1_reg[969 ] <= 8'h00;
memory1_reg[970 ] <= 8'h00;
memory1_reg[971 ] <= 8'h00;
memory1_reg[972 ] <= 8'h00;
memory1_reg[973 ] <= 8'h00;
memory1_reg[974 ] <= 8'h00;
memory1_reg[975 ] <= 8'h00;
memory1_reg[976 ] <= 8'h00;
memory1_reg[977 ] <= 8'h00;
memory1_reg[978 ] <= 8'h00;
memory1_reg[979 ] <= 8'h00;
memory1_reg[980 ] <= 8'h00;
memory1_reg[981 ] <= 8'h00;
memory1_reg[982 ] <= 8'h00;
memory1_reg[983 ] <= 8'h00;
memory1_reg[984 ] <= 8'h00;
memory1_reg[985 ] <= 8'h00;
memory1_reg[986 ] <= 8'h00;
memory1_reg[987 ] <= 8'h00;
memory1_reg[988 ] <= 8'h00;
memory1_reg[989 ] <= 8'h00;
memory1_reg[990 ] <= 8'h00;
memory1_reg[991 ] <= 8'h00;
memory1_reg[992 ] <= 8'h00;
memory1_reg[993 ] <= 8'h00;
memory1_reg[994 ] <= 8'h00;
memory1_reg[995 ] <= 8'h00;
memory1_reg[996 ] <= 8'h00;
memory1_reg[997 ] <= 8'h00;
memory1_reg[998 ] <= 8'h00;
memory1_reg[999 ] <= 8'h00;
memory1_reg[1000] <= 8'h00;
memory1_reg[1001] <= 8'h00;
memory1_reg[1002] <= 8'h00;
memory1_reg[1003] <= 8'h00;
memory1_reg[1004] <= 8'h00;
memory1_reg[1005] <= 8'h00;
memory1_reg[1006] <= 8'h00;
memory1_reg[1007] <= 8'h00;
memory1_reg[1008] <= 8'h00;
memory1_reg[1009] <= 8'h00;
memory1_reg[1010] <= 8'h00;
memory1_reg[1011] <= 8'h00;
memory1_reg[1012] <= 8'h00;
memory1_reg[1013] <= 8'h00;
memory1_reg[1014] <= 8'h00;
memory1_reg[1015] <= 8'h00;
memory1_reg[1016] <= 8'h00;
memory1_reg[1017] <= 8'h00;
memory1_reg[1018] <= 8'h00;
memory1_reg[1019] <= 8'h00;
memory1_reg[1020] <= 8'h00;
memory1_reg[1021] <= 8'h00;
memory1_reg[1022] <= 8'h00;
memory1_reg[1023] <= 8'h00;

// Memory 2

memory2_reg[0   ] <= 8'h00;
memory2_reg[1   ] <= 8'h08;
memory2_reg[2   ] <= 8'h09;
memory2_reg[3   ] <= 8'h08;
memory2_reg[4   ] <= 8'h00;
memory2_reg[5   ] <= 8'h09;
memory2_reg[6   ] <= 8'h0B;
memory2_reg[7   ] <= 8'h08;
memory2_reg[8   ] <= 8'h0B;
memory2_reg[9   ] <= 8'h00;
memory2_reg[10  ] <= 8'h00;
memory2_reg[11  ] <= 8'h08;
memory2_reg[12  ] <= 8'h09;
memory2_reg[13  ] <= 8'h00;
memory2_reg[14  ] <= 8'h09;
memory2_reg[15  ] <= 8'h0B;
memory2_reg[16  ] <= 8'h0B;
memory2_reg[17  ] <= 8'h00;
memory2_reg[18  ] <= 8'h00;
memory2_reg[19  ] <= 8'h08;
memory2_reg[20  ] <= 8'h09;
memory2_reg[21  ] <= 8'h08;
memory2_reg[22  ] <= 8'h00;
memory2_reg[23  ] <= 8'h09;
memory2_reg[24  ] <= 8'h0B;
memory2_reg[25  ] <= 8'h08;
memory2_reg[26  ] <= 8'h0B;
memory2_reg[27  ] <= 8'h00;
memory2_reg[28  ] <= 8'h00;
memory2_reg[29  ] <= 8'h08;
memory2_reg[30  ] <= 8'h09;
memory2_reg[31  ] <= 8'h00;
memory2_reg[32  ] <= 8'h09;
memory2_reg[33  ] <= 8'h0B;
memory2_reg[34  ] <= 8'h0B;
memory2_reg[35  ] <= 8'h00;
memory2_reg[36  ] <= 8'h00;
memory2_reg[37  ] <= 8'h08;
memory2_reg[38  ] <= 8'h09;
memory2_reg[39  ] <= 8'h08;
memory2_reg[40  ] <= 8'h00;
memory2_reg[41  ] <= 8'h09;
memory2_reg[42  ] <= 8'h0B;
memory2_reg[43  ] <= 8'h08;
memory2_reg[44  ] <= 8'h0B;
memory2_reg[45  ] <= 8'h00;
memory2_reg[46  ] <= 8'h00;
memory2_reg[47  ] <= 8'h08;
memory2_reg[48  ] <= 8'h09;
memory2_reg[49  ] <= 8'h00;
memory2_reg[50  ] <= 8'h09;
memory2_reg[51  ] <= 8'h0B;
memory2_reg[52  ] <= 8'h0B;
memory2_reg[53  ] <= 8'h00;
memory2_reg[54  ] <= 8'h00;
memory2_reg[55  ] <= 8'h00;
memory2_reg[56  ] <= 8'h00;
memory2_reg[57  ] <= 8'h08;
memory2_reg[58  ] <= 8'h09;
memory2_reg[59  ] <= 8'h08;
memory2_reg[60  ] <= 8'h00;
memory2_reg[61  ] <= 8'h09;
memory2_reg[62  ] <= 8'h0B;
memory2_reg[63  ] <= 8'h08;
memory2_reg[64  ] <= 8'h0B;
memory2_reg[65  ] <= 8'h00;
memory2_reg[66  ] <= 8'h00;
memory2_reg[67  ] <= 8'h08;
memory2_reg[68  ] <= 8'h09;
memory2_reg[69  ] <= 8'h00;
memory2_reg[70  ] <= 8'h09;
memory2_reg[71  ] <= 8'h0B;
memory2_reg[72  ] <= 8'h0B;
memory2_reg[73  ] <= 8'h00;
memory2_reg[74  ] <= 8'h00;
memory2_reg[75  ] <= 8'h08;
memory2_reg[76  ] <= 8'h09;
memory2_reg[77  ] <= 8'h08;
memory2_reg[78  ] <= 8'h00;
memory2_reg[79  ] <= 8'h09;
memory2_reg[80  ] <= 8'h0B;
memory2_reg[81  ] <= 8'h08;
memory2_reg[82  ] <= 8'h0B;
memory2_reg[83  ] <= 8'h00;
memory2_reg[84  ] <= 8'h00;
memory2_reg[85  ] <= 8'h08;
memory2_reg[86  ] <= 8'h09;
memory2_reg[87  ] <= 8'h00;
memory2_reg[88  ] <= 8'h09;
memory2_reg[89  ] <= 8'h0B;
memory2_reg[90  ] <= 8'h0B;
memory2_reg[91  ] <= 8'h00;
memory2_reg[92  ] <= 8'h00;
memory2_reg[93  ] <= 8'h08;
memory2_reg[94  ] <= 8'h09;
memory2_reg[95  ] <= 8'h08;
memory2_reg[96  ] <= 8'h00;
memory2_reg[97  ] <= 8'h09;
memory2_reg[98  ] <= 8'h0B;
memory2_reg[99  ] <= 8'h08;
memory2_reg[100 ] <= 8'h0B;
memory2_reg[101 ] <= 8'h00;
memory2_reg[102 ] <= 8'h00;
memory2_reg[103 ] <= 8'h08;
memory2_reg[104 ] <= 8'h09;
memory2_reg[105 ] <= 8'h00;
memory2_reg[106 ] <= 8'h09;
memory2_reg[107 ] <= 8'h0B;
memory2_reg[108 ] <= 8'h0B;
memory2_reg[109 ] <= 8'h00;
memory2_reg[110 ] <= 8'h00;
memory2_reg[111 ] <= 8'h00;
memory2_reg[112 ] <= 8'h00;
memory2_reg[113 ] <= 8'h08;
memory2_reg[114 ] <= 8'h09;
memory2_reg[115 ] <= 8'h08;
memory2_reg[116 ] <= 8'h00;
memory2_reg[117 ] <= 8'h09;
memory2_reg[118 ] <= 8'h0B;
memory2_reg[119 ] <= 8'h08;
memory2_reg[120 ] <= 8'h0B;
memory2_reg[121 ] <= 8'h00;
memory2_reg[122 ] <= 8'h00;
memory2_reg[123 ] <= 8'h08;
memory2_reg[124 ] <= 8'h09;
memory2_reg[125 ] <= 8'h00;
memory2_reg[126 ] <= 8'h09;
memory2_reg[127 ] <= 8'h0B;
memory2_reg[128 ] <= 8'h0B;
memory2_reg[129 ] <= 8'h00;
memory2_reg[130 ] <= 8'h00;
memory2_reg[131 ] <= 8'h08;
memory2_reg[132 ] <= 8'h09;
memory2_reg[133 ] <= 8'h08;
memory2_reg[134 ] <= 8'h00;
memory2_reg[135 ] <= 8'h09;
memory2_reg[136 ] <= 8'h0B;
memory2_reg[137 ] <= 8'h08;
memory2_reg[138 ] <= 8'h0B;
memory2_reg[139 ] <= 8'h00;
memory2_reg[140 ] <= 8'h00;
memory2_reg[141 ] <= 8'h08;
memory2_reg[142 ] <= 8'h09;
memory2_reg[143 ] <= 8'h00;
memory2_reg[144 ] <= 8'h09;
memory2_reg[145 ] <= 8'h0B;
memory2_reg[146 ] <= 8'h0B;
memory2_reg[147 ] <= 8'h00;
memory2_reg[148 ] <= 8'h00;
memory2_reg[149 ] <= 8'h08;
memory2_reg[150 ] <= 8'h09;
memory2_reg[151 ] <= 8'h08;
memory2_reg[152 ] <= 8'h00;
memory2_reg[153 ] <= 8'h09;
memory2_reg[154 ] <= 8'h0B;
memory2_reg[155 ] <= 8'h08;
memory2_reg[156 ] <= 8'h0B;
memory2_reg[157 ] <= 8'h00;
memory2_reg[158 ] <= 8'h00;
memory2_reg[159 ] <= 8'h08;
memory2_reg[160 ] <= 8'h09;
memory2_reg[161 ] <= 8'h00;
memory2_reg[162 ] <= 8'h09;
memory2_reg[163 ] <= 8'h0B;
memory2_reg[164 ] <= 8'h0B;
memory2_reg[165 ] <= 8'h00;
memory2_reg[166 ] <= 8'h00;
memory2_reg[167 ] <= 8'h00;
memory2_reg[168 ] <= 8'h00;
memory2_reg[169 ] <= 8'h0A;
memory2_reg[170 ] <= 8'h09;
memory2_reg[171 ] <= 8'h00;
memory2_reg[172 ] <= 8'h0A;
memory2_reg[173 ] <= 8'h09;
memory2_reg[174 ] <= 8'h00;
memory2_reg[175 ] <= 8'h0A;
memory2_reg[176 ] <= 8'h09;
memory2_reg[177 ] <= 8'h08;
memory2_reg[178 ] <= 8'h00;
memory2_reg[179 ] <= 8'h0A;
memory2_reg[180 ] <= 8'h09;
memory2_reg[181 ] <= 8'h00;
memory2_reg[182 ] <= 8'h0A;
memory2_reg[183 ] <= 8'h09;
memory2_reg[184 ] <= 8'h00;
memory2_reg[185 ] <= 8'h0A;
memory2_reg[186 ] <= 8'h09;
memory2_reg[187 ] <= 8'h08;
memory2_reg[188 ] <= 8'h00;
memory2_reg[189 ] <= 8'h0A;
memory2_reg[190 ] <= 8'h09;
memory2_reg[191 ] <= 8'h00;
memory2_reg[192 ] <= 8'h0A;
memory2_reg[193 ] <= 8'h09;
memory2_reg[194 ] <= 8'h00;
memory2_reg[195 ] <= 8'h0A;
memory2_reg[196 ] <= 8'h09;
memory2_reg[197 ] <= 8'h08;
memory2_reg[198 ] <= 8'h00;
memory2_reg[199 ] <= 8'h00;
memory2_reg[200 ] <= 8'h00;
memory2_reg[201 ] <= 8'h00;
memory2_reg[202 ] <= 8'h00;
memory2_reg[203 ] <= 8'h00;
memory2_reg[204 ] <= 8'h00;
memory2_reg[205 ] <= 8'h00;
memory2_reg[206 ] <= 8'h00;
memory2_reg[207 ] <= 8'h00;
memory2_reg[208 ] <= 8'h00;
memory2_reg[209 ] <= 8'h00;
memory2_reg[210 ] <= 8'h00;
memory2_reg[211 ] <= 8'h00;
memory2_reg[212 ] <= 8'h00;
memory2_reg[213 ] <= 8'h00;
memory2_reg[214 ] <= 8'h00;
memory2_reg[215 ] <= 8'h00;
memory2_reg[216 ] <= 8'h00;
memory2_reg[217 ] <= 8'h00;
memory2_reg[218 ] <= 8'h00;
memory2_reg[219 ] <= 8'h00;
memory2_reg[220 ] <= 8'h00;
memory2_reg[221 ] <= 8'h00;
memory2_reg[222 ] <= 8'h00;
memory2_reg[223 ] <= 8'h00;
memory2_reg[224 ] <= 8'h00;
memory2_reg[225 ] <= 8'h00;
memory2_reg[226 ] <= 8'h00;
memory2_reg[227 ] <= 8'h00;
memory2_reg[228 ] <= 8'h00;
memory2_reg[229 ] <= 8'h00;
memory2_reg[230 ] <= 8'h00;
memory2_reg[231 ] <= 8'h00;
memory2_reg[232 ] <= 8'h00;
memory2_reg[233 ] <= 8'h00;
memory2_reg[234 ] <= 8'h00;
memory2_reg[235 ] <= 8'h00;
memory2_reg[236 ] <= 8'h00;
memory2_reg[237 ] <= 8'h00;
memory2_reg[238 ] <= 8'h00;
memory2_reg[239 ] <= 8'h00;
memory2_reg[240 ] <= 8'h00;
memory2_reg[241 ] <= 8'h00;
memory2_reg[242 ] <= 8'h00;
memory2_reg[243 ] <= 8'h00;
memory2_reg[244 ] <= 8'h00;
memory2_reg[245 ] <= 8'h00;
memory2_reg[246 ] <= 8'h00;
memory2_reg[247 ] <= 8'h00;
memory2_reg[248 ] <= 8'h00;
memory2_reg[249 ] <= 8'h00;
memory2_reg[250 ] <= 8'h00;
memory2_reg[251 ] <= 8'h00;
memory2_reg[252 ] <= 8'h00;
memory2_reg[253 ] <= 8'h00;
memory2_reg[254 ] <= 8'h00;
memory2_reg[255 ] <= 8'h00;
memory2_reg[256 ] <= 8'h08;
memory2_reg[257 ] <= 8'h0A;
memory2_reg[258 ] <= 8'h09;
memory2_reg[259 ] <= 8'h0A;
memory2_reg[260 ] <= 8'h09;
memory2_reg[261 ] <= 8'h0A;
memory2_reg[262 ] <= 8'h09;
memory2_reg[263 ] <= 8'h08;
memory2_reg[264 ] <= 8'h0A;
memory2_reg[265 ] <= 8'h09;
memory2_reg[266 ] <= 8'h0A;
memory2_reg[267 ] <= 8'h09;
memory2_reg[268 ] <= 8'h0A;
memory2_reg[269 ] <= 8'h09;
memory2_reg[270 ] <= 8'h08;
memory2_reg[271 ] <= 8'h0A;
memory2_reg[272 ] <= 8'h09;
memory2_reg[273 ] <= 8'h0A;
memory2_reg[274 ] <= 8'h09;
memory2_reg[275 ] <= 8'h0A;
memory2_reg[276 ] <= 8'h09;
memory2_reg[277 ] <= 8'h08;
memory2_reg[278 ] <= 8'h0A;
memory2_reg[279 ] <= 8'h09;
memory2_reg[280 ] <= 8'h0A;
memory2_reg[281 ] <= 8'h09;
memory2_reg[282 ] <= 8'h0A;
memory2_reg[283 ] <= 8'h09;
memory2_reg[284 ] <= 8'h08;
memory2_reg[285 ] <= 8'h0A;
memory2_reg[286 ] <= 8'h09;
memory2_reg[287 ] <= 8'h0A;
memory2_reg[288 ] <= 8'h09;
memory2_reg[289 ] <= 8'h0A;
memory2_reg[290 ] <= 8'h09;
memory2_reg[291 ] <= 8'h08;
memory2_reg[292 ] <= 8'h0A;
memory2_reg[293 ] <= 8'h09;
memory2_reg[294 ] <= 8'h0A;
memory2_reg[295 ] <= 8'h09;
memory2_reg[296 ] <= 8'h0A;
memory2_reg[297 ] <= 8'h09;
memory2_reg[298 ] <= 8'h08;
memory2_reg[299 ] <= 8'h0A;
memory2_reg[300 ] <= 8'h09;
memory2_reg[301 ] <= 8'h0A;
memory2_reg[302 ] <= 8'h09;
memory2_reg[303 ] <= 8'h0A;
memory2_reg[304 ] <= 8'h09;
memory2_reg[305 ] <= 8'h08;
memory2_reg[306 ] <= 8'h0A;
memory2_reg[307 ] <= 8'h09;
memory2_reg[308 ] <= 8'h0A;
memory2_reg[309 ] <= 8'h09;
memory2_reg[310 ] <= 8'h0A;
memory2_reg[311 ] <= 8'h09;
memory2_reg[312 ] <= 8'h08;
memory2_reg[313 ] <= 8'h0A;
memory2_reg[314 ] <= 8'h09;
memory2_reg[315 ] <= 8'h0A;
memory2_reg[316 ] <= 8'h09;
memory2_reg[317 ] <= 8'h0A;
memory2_reg[318 ] <= 8'h09;
memory2_reg[319 ] <= 8'h08;
memory2_reg[320 ] <= 8'h08;
memory2_reg[321 ] <= 8'h08;
memory2_reg[322 ] <= 8'h00;
memory2_reg[323 ] <= 8'h08;
memory2_reg[324 ] <= 8'h00;
memory2_reg[325 ] <= 8'h08;
memory2_reg[326 ] <= 8'h00;
memory2_reg[327 ] <= 8'h08;
memory2_reg[328 ] <= 8'h08;
memory2_reg[329 ] <= 8'h08;
memory2_reg[330 ] <= 8'h00;
memory2_reg[331 ] <= 8'h08;
memory2_reg[332 ] <= 8'h00;
memory2_reg[333 ] <= 8'h08;
memory2_reg[334 ] <= 8'h00;
memory2_reg[335 ] <= 8'h08;
memory2_reg[336 ] <= 8'h08;
memory2_reg[337 ] <= 8'h08;
memory2_reg[338 ] <= 8'h00;
memory2_reg[339 ] <= 8'h08;
memory2_reg[340 ] <= 8'h00;
memory2_reg[341 ] <= 8'h08;
memory2_reg[342 ] <= 8'h00;
memory2_reg[343 ] <= 8'h08;
memory2_reg[344 ] <= 8'h08;
memory2_reg[345 ] <= 8'h08;
memory2_reg[346 ] <= 8'h0B;
memory2_reg[347 ] <= 8'h0B;
memory2_reg[348 ] <= 8'h08;
memory2_reg[349 ] <= 8'h00;
memory2_reg[350 ] <= 8'h00;
memory2_reg[351 ] <= 8'h00;
memory2_reg[352 ] <= 8'h08;
memory2_reg[353 ] <= 8'h00;
memory2_reg[354 ] <= 8'h00;
memory2_reg[355 ] <= 8'h00;
memory2_reg[356 ] <= 8'h08;
memory2_reg[357 ] <= 8'h00;
memory2_reg[358 ] <= 8'h00;
memory2_reg[359 ] <= 8'h00;
memory2_reg[360 ] <= 8'h00;
memory2_reg[361 ] <= 8'h00;
memory2_reg[362 ] <= 8'h00;
memory2_reg[363 ] <= 8'h00;
memory2_reg[364 ] <= 8'h00;
memory2_reg[365 ] <= 8'h00;
memory2_reg[366 ] <= 8'h00;
memory2_reg[367 ] <= 8'h00;
memory2_reg[368 ] <= 8'h08;
memory2_reg[369 ] <= 8'h08;
memory2_reg[370 ] <= 8'h00;
memory2_reg[371 ] <= 8'h00;
memory2_reg[372 ] <= 8'h08;
memory2_reg[373 ] <= 8'h08;
memory2_reg[374 ] <= 8'h08;
memory2_reg[375 ] <= 8'h08;
memory2_reg[376 ] <= 8'h08;
memory2_reg[377 ] <= 8'h08;
memory2_reg[378 ] <= 8'h08;
memory2_reg[379 ] <= 8'h08;
memory2_reg[380 ] <= 8'h00;
memory2_reg[381 ] <= 8'h08;
memory2_reg[382 ] <= 8'h09;
memory2_reg[383 ] <= 8'h08;
memory2_reg[384 ] <= 8'h08;
memory2_reg[385 ] <= 8'h0A;
memory2_reg[386 ] <= 8'h00;
memory2_reg[387 ] <= 8'h09;
memory2_reg[388 ] <= 8'h00;
memory2_reg[389 ] <= 8'h09;
memory2_reg[390 ] <= 8'h00;
memory2_reg[391 ] <= 8'h09;
memory2_reg[392 ] <= 8'h08;
memory2_reg[393 ] <= 8'h0A;
memory2_reg[394 ] <= 8'h00;
memory2_reg[395 ] <= 8'h09;
memory2_reg[396 ] <= 8'h00;
memory2_reg[397 ] <= 8'h09;
memory2_reg[398 ] <= 8'h00;
memory2_reg[399 ] <= 8'h09;
memory2_reg[400 ] <= 8'h08;
memory2_reg[401 ] <= 8'h0A;
memory2_reg[402 ] <= 8'h00;
memory2_reg[403 ] <= 8'h09;
memory2_reg[404 ] <= 8'h00;
memory2_reg[405 ] <= 8'h09;
memory2_reg[406 ] <= 8'h00;
memory2_reg[407 ] <= 8'h09;
memory2_reg[408 ] <= 8'h08;
memory2_reg[409 ] <= 8'h00;
memory2_reg[410 ] <= 8'h00;
memory2_reg[411 ] <= 8'h00;
memory2_reg[412 ] <= 8'h00;
memory2_reg[413 ] <= 8'h0A;
memory2_reg[414 ] <= 8'h09;
memory2_reg[415 ] <= 8'h08;
memory2_reg[416 ] <= 8'h08;
memory2_reg[417 ] <= 8'h08;
memory2_reg[418 ] <= 8'h09;
memory2_reg[419 ] <= 8'h08;
memory2_reg[420 ] <= 8'h00;
memory2_reg[421 ] <= 8'h0A;
memory2_reg[422 ] <= 8'h09;
memory2_reg[423 ] <= 8'h08;
memory2_reg[424 ] <= 8'h08;
memory2_reg[425 ] <= 8'h08;
memory2_reg[426 ] <= 8'h09;
memory2_reg[427 ] <= 8'h08;
memory2_reg[428 ] <= 8'h00;
memory2_reg[429 ] <= 8'h0A;
memory2_reg[430 ] <= 8'h09;
memory2_reg[431 ] <= 8'h08;
memory2_reg[432 ] <= 8'h08;
memory2_reg[433 ] <= 8'h08;
memory2_reg[434 ] <= 8'h09;
memory2_reg[435 ] <= 8'h08;
memory2_reg[436 ] <= 8'h08;
memory2_reg[437 ] <= 8'h08;
memory2_reg[438 ] <= 8'h09;
memory2_reg[439 ] <= 8'h08;
memory2_reg[440 ] <= 8'h09;
memory2_reg[441 ] <= 8'h08;
memory2_reg[442 ] <= 8'h09;
memory2_reg[443 ] <= 8'h08;
memory2_reg[444 ] <= 8'h08;
memory2_reg[445 ] <= 8'h09;
memory2_reg[446 ] <= 8'h08;
memory2_reg[447 ] <= 8'h09;
memory2_reg[448 ] <= 8'h08;
memory2_reg[449 ] <= 8'h09;
memory2_reg[450 ] <= 8'h08;
memory2_reg[451 ] <= 8'h08;
memory2_reg[452 ] <= 8'h09;
memory2_reg[453 ] <= 8'h08;
memory2_reg[454 ] <= 8'h09;
memory2_reg[455 ] <= 8'h08;
memory2_reg[456 ] <= 8'h09;
memory2_reg[457 ] <= 8'h08;
memory2_reg[458 ] <= 8'h08;
memory2_reg[459 ] <= 8'h0B;
memory2_reg[460 ] <= 8'h0B;
memory2_reg[461 ] <= 8'h0B;
memory2_reg[462 ] <= 8'h0B;
memory2_reg[463 ] <= 8'h0B;
memory2_reg[464 ] <= 8'h08;
memory2_reg[465 ] <= 8'h08;
memory2_reg[466 ] <= 8'h0B;
memory2_reg[467 ] <= 8'h08;
memory2_reg[468 ] <= 8'h08;
memory2_reg[469 ] <= 8'h0B;
memory2_reg[470 ] <= 8'h08;
memory2_reg[471 ] <= 8'h08;
memory2_reg[472 ] <= 8'h0B;
memory2_reg[473 ] <= 8'h00;
memory2_reg[474 ] <= 8'h00;
memory2_reg[475 ] <= 8'h00;
memory2_reg[476 ] <= 8'h00;
memory2_reg[477 ] <= 8'h09;
memory2_reg[478 ] <= 8'h00;
memory2_reg[479 ] <= 8'h09;
memory2_reg[480 ] <= 8'h00;
memory2_reg[481 ] <= 8'h09;
memory2_reg[482 ] <= 8'h00;
memory2_reg[483 ] <= 8'h09;
memory2_reg[484 ] <= 8'h00;
memory2_reg[485 ] <= 8'h09;
memory2_reg[486 ] <= 8'h00;
memory2_reg[487 ] <= 8'h09;
memory2_reg[488 ] <= 8'h00;
memory2_reg[489 ] <= 8'h09;
memory2_reg[490 ] <= 8'h00;
memory2_reg[491 ] <= 8'h09;
memory2_reg[492 ] <= 8'h00;
memory2_reg[493 ] <= 8'h09;
memory2_reg[494 ] <= 8'h00;
memory2_reg[495 ] <= 8'h0A;
memory2_reg[496 ] <= 8'h00;
memory2_reg[497 ] <= 8'h0A;
memory2_reg[498 ] <= 8'h00;
memory2_reg[499 ] <= 8'h0A;
memory2_reg[500 ] <= 8'h00;
memory2_reg[501 ] <= 8'h00;
memory2_reg[502 ] <= 8'h00;
memory2_reg[503 ] <= 8'h00;
memory2_reg[504 ] <= 8'h00;
memory2_reg[505 ] <= 8'h00;
memory2_reg[506 ] <= 8'h00;
memory2_reg[507 ] <= 8'h00;
memory2_reg[508 ] <= 8'h00;
memory2_reg[509 ] <= 8'h00;
memory2_reg[510 ] <= 8'h00;
memory2_reg[511 ] <= 8'h00;
memory2_reg[512 ] <= 8'h00;
memory2_reg[513 ] <= 8'h0A;
memory2_reg[514 ] <= 8'h00;
memory2_reg[515 ] <= 8'h0A;
memory2_reg[516 ] <= 8'h00;
memory2_reg[517 ] <= 8'h0A;
memory2_reg[518 ] <= 8'h00;
memory2_reg[519 ] <= 8'h0A;
memory2_reg[520 ] <= 8'h00;
memory2_reg[521 ] <= 8'h0A;
memory2_reg[522 ] <= 8'h00;
memory2_reg[523 ] <= 8'h0A;
memory2_reg[524 ] <= 8'h00;
memory2_reg[525 ] <= 8'h0A;
memory2_reg[526 ] <= 8'h00;
memory2_reg[527 ] <= 8'h0A;
memory2_reg[528 ] <= 8'h00;
memory2_reg[529 ] <= 8'h0A;
memory2_reg[530 ] <= 8'h00;
memory2_reg[531 ] <= 8'h0B;
memory2_reg[532 ] <= 8'h00;
memory2_reg[533 ] <= 8'h0B;
memory2_reg[534 ] <= 8'h00;
memory2_reg[535 ] <= 8'h0B;
memory2_reg[536 ] <= 8'h08;
memory2_reg[537 ] <= 8'h08;
memory2_reg[538 ] <= 8'h08;
memory2_reg[539 ] <= 8'h08;
memory2_reg[540 ] <= 8'h08;
memory2_reg[541 ] <= 8'h08;
memory2_reg[542 ] <= 8'h08;
memory2_reg[543 ] <= 8'h00;
memory2_reg[544 ] <= 8'h08;
memory2_reg[545 ] <= 8'h09;
memory2_reg[546 ] <= 8'h09;
memory2_reg[547 ] <= 8'h09;
memory2_reg[548 ] <= 8'h09;
memory2_reg[549 ] <= 8'h0B;
memory2_reg[550 ] <= 8'h00;
memory2_reg[551 ] <= 8'h00;
memory2_reg[552 ] <= 8'h0B;
memory2_reg[553 ] <= 8'h0B;
memory2_reg[554 ] <= 8'h0B;
memory2_reg[555 ] <= 8'h0B;
memory2_reg[556 ] <= 8'h09;
memory2_reg[557 ] <= 8'h0B;
memory2_reg[558 ] <= 8'h0B;
memory2_reg[559 ] <= 8'h09;
memory2_reg[560 ] <= 8'h0B;
memory2_reg[561 ] <= 8'h09;
memory2_reg[562 ] <= 8'h0B;
memory2_reg[563 ] <= 8'h09;
memory2_reg[564 ] <= 8'h08;
memory2_reg[565 ] <= 8'h09;
memory2_reg[566 ] <= 8'h09;
memory2_reg[567 ] <= 8'h0B;
memory2_reg[568 ] <= 8'h09;
memory2_reg[569 ] <= 8'h0B;
memory2_reg[570 ] <= 8'h09;
memory2_reg[571 ] <= 8'h0B;
memory2_reg[572 ] <= 8'h09;
memory2_reg[573 ] <= 8'h08;
memory2_reg[574 ] <= 8'h09;
memory2_reg[575 ] <= 8'h09;
memory2_reg[576 ] <= 8'h0B;
memory2_reg[577 ] <= 8'h09;
memory2_reg[578 ] <= 8'h0B;
memory2_reg[579 ] <= 8'h09;
memory2_reg[580 ] <= 8'h09;
memory2_reg[581 ] <= 8'h0B;
memory2_reg[582 ] <= 8'h09;
memory2_reg[583 ] <= 8'h09;
memory2_reg[584 ] <= 8'h0B;
memory2_reg[585 ] <= 8'h09;
memory2_reg[586 ] <= 8'h0B;
memory2_reg[587 ] <= 8'h08;
memory2_reg[588 ] <= 8'h09;
memory2_reg[589 ] <= 8'h09;
memory2_reg[590 ] <= 8'h0B;
memory2_reg[591 ] <= 8'h09;
memory2_reg[592 ] <= 8'h09;
memory2_reg[593 ] <= 8'h0B;
memory2_reg[594 ] <= 8'h09;
memory2_reg[595 ] <= 8'h0B;
memory2_reg[596 ] <= 8'h08;
memory2_reg[597 ] <= 8'h0A;
memory2_reg[598 ] <= 8'h08;
memory2_reg[599 ] <= 8'h0A;
memory2_reg[600 ] <= 8'h08;
memory2_reg[601 ] <= 8'h09;
memory2_reg[602 ] <= 8'h09;
memory2_reg[603 ] <= 8'h09;
memory2_reg[604 ] <= 8'h09;
memory2_reg[605 ] <= 8'h09;
memory2_reg[606 ] <= 8'h09;
memory2_reg[607 ] <= 8'h0B;
memory2_reg[608 ] <= 8'h0A;
memory2_reg[609 ] <= 8'h09;
memory2_reg[610 ] <= 8'h08;
memory2_reg[611 ] <= 8'h09;
memory2_reg[612 ] <= 8'h0B;
memory2_reg[613 ] <= 8'h09;
memory2_reg[614 ] <= 8'h0A;
memory2_reg[615 ] <= 8'h0A;
memory2_reg[616 ] <= 8'h09;
memory2_reg[617 ] <= 8'h08;
memory2_reg[618 ] <= 8'h09;
memory2_reg[619 ] <= 8'h0B;
memory2_reg[620 ] <= 8'h09;
memory2_reg[621 ] <= 8'h0A;
memory2_reg[622 ] <= 8'h0B;
memory2_reg[623 ] <= 8'h0A;
memory2_reg[624 ] <= 8'h09;
memory2_reg[625 ] <= 8'h08;
memory2_reg[626 ] <= 8'h09;
memory2_reg[627 ] <= 8'h0B;
memory2_reg[628 ] <= 8'h09;
memory2_reg[629 ] <= 8'h0A;
memory2_reg[630 ] <= 8'h00;
memory2_reg[631 ] <= 8'h00;
memory2_reg[632 ] <= 8'h08;
memory2_reg[633 ] <= 8'h0A;
memory2_reg[634 ] <= 8'h08;
memory2_reg[635 ] <= 8'h0A;
memory2_reg[636 ] <= 8'h0A;
memory2_reg[637 ] <= 8'h09;
memory2_reg[638 ] <= 8'h08;
memory2_reg[639 ] <= 8'h09;
memory2_reg[640 ] <= 8'h0A;
memory2_reg[641 ] <= 8'h0A;
memory2_reg[642 ] <= 8'h09;
memory2_reg[643 ] <= 8'h08;
memory2_reg[644 ] <= 8'h09;
memory2_reg[645 ] <= 8'h0A;
memory2_reg[646 ] <= 8'h0B;
memory2_reg[647 ] <= 8'h0A;
memory2_reg[648 ] <= 8'h09;
memory2_reg[649 ] <= 8'h08;
memory2_reg[650 ] <= 8'h09;
memory2_reg[651 ] <= 8'h0A;
memory2_reg[652 ] <= 8'h08;
memory2_reg[653 ] <= 8'h0A;
memory2_reg[654 ] <= 8'h08;
memory2_reg[655 ] <= 8'h0A;
memory2_reg[656 ] <= 8'h08;
memory2_reg[657 ] <= 8'h09;
memory2_reg[658 ] <= 8'h09;
memory2_reg[659 ] <= 8'h09;
memory2_reg[660 ] <= 8'h09;
memory2_reg[661 ] <= 8'h09;
memory2_reg[662 ] <= 8'h09;
memory2_reg[663 ] <= 8'h0B;
memory2_reg[664 ] <= 8'h08;
memory2_reg[665 ] <= 8'h0A;
memory2_reg[666 ] <= 8'h09;
memory2_reg[667 ] <= 8'h08;
memory2_reg[668 ] <= 8'h09;
memory2_reg[669 ] <= 8'h0B;
memory2_reg[670 ] <= 8'h09;
memory2_reg[671 ] <= 8'h0A;
memory2_reg[672 ] <= 8'h0A;
memory2_reg[673 ] <= 8'h09;
memory2_reg[674 ] <= 8'h08;
memory2_reg[675 ] <= 8'h09;
memory2_reg[676 ] <= 8'h0B;
memory2_reg[677 ] <= 8'h09;
memory2_reg[678 ] <= 8'h0A;
memory2_reg[679 ] <= 8'h0B;
memory2_reg[680 ] <= 8'h0A;
memory2_reg[681 ] <= 8'h09;
memory2_reg[682 ] <= 8'h08;
memory2_reg[683 ] <= 8'h09;
memory2_reg[684 ] <= 8'h0B;
memory2_reg[685 ] <= 8'h09;
memory2_reg[686 ] <= 8'h0A;
memory2_reg[687 ] <= 8'h00;
memory2_reg[688 ] <= 8'h08;
memory2_reg[689 ] <= 8'h09;
memory2_reg[690 ] <= 8'h09;
memory2_reg[691 ] <= 8'h09;
memory2_reg[692 ] <= 8'h09;
memory2_reg[693 ] <= 8'h09;
memory2_reg[694 ] <= 8'h09;
memory2_reg[695 ] <= 8'h0B;
memory2_reg[696 ] <= 8'h00;
memory2_reg[697 ] <= 8'h08;
memory2_reg[698 ] <= 8'h08;
memory2_reg[699 ] <= 8'h00;
memory2_reg[700 ] <= 8'h00;
memory2_reg[701 ] <= 8'h08;
memory2_reg[702 ] <= 8'h08;
memory2_reg[703 ] <= 8'h00;
memory2_reg[704 ] <= 8'h00;
memory2_reg[705 ] <= 8'h08;
memory2_reg[706 ] <= 8'h09;
memory2_reg[707 ] <= 8'h08;
memory2_reg[708 ] <= 8'h00;
memory2_reg[709 ] <= 8'h00;
memory2_reg[710 ] <= 8'h00;
memory2_reg[711 ] <= 8'h00;
memory2_reg[712 ] <= 8'h00;
memory2_reg[713 ] <= 8'h00;
memory2_reg[714 ] <= 8'h00;
memory2_reg[715 ] <= 8'h00;
memory2_reg[716 ] <= 8'h00;
memory2_reg[717 ] <= 8'h00;
memory2_reg[718 ] <= 8'h00;
memory2_reg[719 ] <= 8'h00;
memory2_reg[720 ] <= 8'h00;
memory2_reg[721 ] <= 8'h00;
memory2_reg[722 ] <= 8'h00;
memory2_reg[723 ] <= 8'h00;
memory2_reg[724 ] <= 8'h00;
memory2_reg[725 ] <= 8'h00;
memory2_reg[726 ] <= 8'h00;
memory2_reg[727 ] <= 8'h00;
memory2_reg[728 ] <= 8'h00;
memory2_reg[729 ] <= 8'h00;
memory2_reg[730 ] <= 8'h00;
memory2_reg[731 ] <= 8'h00;
memory2_reg[732 ] <= 8'h00;
memory2_reg[733 ] <= 8'h00;
memory2_reg[734 ] <= 8'h00;
memory2_reg[735 ] <= 8'h00;
memory2_reg[736 ] <= 8'h00;
memory2_reg[737 ] <= 8'h00;
memory2_reg[738 ] <= 8'h00;
memory2_reg[739 ] <= 8'h00;
memory2_reg[740 ] <= 8'h00;
memory2_reg[741 ] <= 8'h00;
memory2_reg[742 ] <= 8'h00;
memory2_reg[743 ] <= 8'h00;
memory2_reg[744 ] <= 8'h00;
memory2_reg[745 ] <= 8'h00;
memory2_reg[746 ] <= 8'h00;
memory2_reg[747 ] <= 8'h00;
memory2_reg[748 ] <= 8'h00;
memory2_reg[749 ] <= 8'h00;
memory2_reg[750 ] <= 8'h00;
memory2_reg[751 ] <= 8'h00;
memory2_reg[752 ] <= 8'h00;
memory2_reg[753 ] <= 8'h00;
memory2_reg[754 ] <= 8'h00;
memory2_reg[755 ] <= 8'h00;
memory2_reg[756 ] <= 8'h00;
memory2_reg[757 ] <= 8'h00;
memory2_reg[758 ] <= 8'h00;
memory2_reg[759 ] <= 8'h00;
memory2_reg[760 ] <= 8'h00;
memory2_reg[761 ] <= 8'h00;
memory2_reg[762 ] <= 8'h00;
memory2_reg[763 ] <= 8'h00;
memory2_reg[764 ] <= 8'h00;
memory2_reg[765 ] <= 8'h00;
memory2_reg[766 ] <= 8'h00;
memory2_reg[767 ] <= 8'h00;
memory2_reg[768 ] <= 8'h00;
memory2_reg[769 ] <= 8'h00;
memory2_reg[770 ] <= 8'h00;
memory2_reg[771 ] <= 8'h00;
memory2_reg[772 ] <= 8'h00;
memory2_reg[773 ] <= 8'h00;
memory2_reg[774 ] <= 8'h00;
memory2_reg[775 ] <= 8'h00;
memory2_reg[776 ] <= 8'h00;
memory2_reg[777 ] <= 8'h00;
memory2_reg[778 ] <= 8'h00;
memory2_reg[779 ] <= 8'h00;
memory2_reg[780 ] <= 8'h00;
memory2_reg[781 ] <= 8'h00;
memory2_reg[782 ] <= 8'h00;
memory2_reg[783 ] <= 8'h00;
memory2_reg[784 ] <= 8'h00;
memory2_reg[785 ] <= 8'h00;
memory2_reg[786 ] <= 8'h00;
memory2_reg[787 ] <= 8'h00;
memory2_reg[788 ] <= 8'h00;
memory2_reg[789 ] <= 8'h00;
memory2_reg[790 ] <= 8'h00;
memory2_reg[791 ] <= 8'h00;
memory2_reg[792 ] <= 8'h00;
memory2_reg[793 ] <= 8'h00;
memory2_reg[794 ] <= 8'h00;
memory2_reg[795 ] <= 8'h00;
memory2_reg[796 ] <= 8'h00;
memory2_reg[797 ] <= 8'h00;
memory2_reg[798 ] <= 8'h00;
memory2_reg[799 ] <= 8'h00;
memory2_reg[800 ] <= 8'h00;
memory2_reg[801 ] <= 8'h00;
memory2_reg[802 ] <= 8'h00;
memory2_reg[803 ] <= 8'h00;
memory2_reg[804 ] <= 8'h00;
memory2_reg[805 ] <= 8'h00;
memory2_reg[806 ] <= 8'h00;
memory2_reg[807 ] <= 8'h00;
memory2_reg[808 ] <= 8'h00;
memory2_reg[809 ] <= 8'h00;
memory2_reg[810 ] <= 8'h00;
memory2_reg[811 ] <= 8'h00;
memory2_reg[812 ] <= 8'h00;
memory2_reg[813 ] <= 8'h00;
memory2_reg[814 ] <= 8'h00;
memory2_reg[815 ] <= 8'h00;
memory2_reg[816 ] <= 8'h00;
memory2_reg[817 ] <= 8'h00;
memory2_reg[818 ] <= 8'h00;
memory2_reg[819 ] <= 8'h00;
memory2_reg[820 ] <= 8'h00;
memory2_reg[821 ] <= 8'h00;
memory2_reg[822 ] <= 8'h00;
memory2_reg[823 ] <= 8'h00;
memory2_reg[824 ] <= 8'h00;
memory2_reg[825 ] <= 8'h00;
memory2_reg[826 ] <= 8'h00;
memory2_reg[827 ] <= 8'h00;
memory2_reg[828 ] <= 8'h00;
memory2_reg[829 ] <= 8'h00;
memory2_reg[830 ] <= 8'h00;
memory2_reg[831 ] <= 8'h00;
memory2_reg[832 ] <= 8'h00;
memory2_reg[833 ] <= 8'h00;
memory2_reg[834 ] <= 8'h00;
memory2_reg[835 ] <= 8'h00;
memory2_reg[836 ] <= 8'h00;
memory2_reg[837 ] <= 8'h00;
memory2_reg[838 ] <= 8'h00;
memory2_reg[839 ] <= 8'h00;
memory2_reg[840 ] <= 8'h00;
memory2_reg[841 ] <= 8'h00;
memory2_reg[842 ] <= 8'h00;
memory2_reg[843 ] <= 8'h00;
memory2_reg[844 ] <= 8'h00;
memory2_reg[845 ] <= 8'h00;
memory2_reg[846 ] <= 8'h00;
memory2_reg[847 ] <= 8'h00;
memory2_reg[848 ] <= 8'h00;
memory2_reg[849 ] <= 8'h00;
memory2_reg[850 ] <= 8'h00;
memory2_reg[851 ] <= 8'h00;
memory2_reg[852 ] <= 8'h00;
memory2_reg[853 ] <= 8'h00;
memory2_reg[854 ] <= 8'h00;
memory2_reg[855 ] <= 8'h00;
memory2_reg[856 ] <= 8'h00;
memory2_reg[857 ] <= 8'h00;
memory2_reg[858 ] <= 8'h00;
memory2_reg[859 ] <= 8'h00;
memory2_reg[860 ] <= 8'h00;
memory2_reg[861 ] <= 8'h00;
memory2_reg[862 ] <= 8'h00;
memory2_reg[863 ] <= 8'h00;
memory2_reg[864 ] <= 8'h00;
memory2_reg[865 ] <= 8'h00;
memory2_reg[866 ] <= 8'h00;
memory2_reg[867 ] <= 8'h00;
memory2_reg[868 ] <= 8'h00;
memory2_reg[869 ] <= 8'h00;
memory2_reg[870 ] <= 8'h00;
memory2_reg[871 ] <= 8'h00;
memory2_reg[872 ] <= 8'h00;
memory2_reg[873 ] <= 8'h00;
memory2_reg[874 ] <= 8'h00;
memory2_reg[875 ] <= 8'h00;
memory2_reg[876 ] <= 8'h00;
memory2_reg[877 ] <= 8'h00;
memory2_reg[878 ] <= 8'h00;
memory2_reg[879 ] <= 8'h00;
memory2_reg[880 ] <= 8'h00;
memory2_reg[881 ] <= 8'h00;
memory2_reg[882 ] <= 8'h00;
memory2_reg[883 ] <= 8'h00;
memory2_reg[884 ] <= 8'h00;
memory2_reg[885 ] <= 8'h00;
memory2_reg[886 ] <= 8'h00;
memory2_reg[887 ] <= 8'h00;
memory2_reg[888 ] <= 8'h00;
memory2_reg[889 ] <= 8'h00;
memory2_reg[890 ] <= 8'h00;
memory2_reg[891 ] <= 8'h00;
memory2_reg[892 ] <= 8'h00;
memory2_reg[893 ] <= 8'h00;
memory2_reg[894 ] <= 8'h00;
memory2_reg[895 ] <= 8'h00;
memory2_reg[896 ] <= 8'h00;
memory2_reg[897 ] <= 8'h00;
memory2_reg[898 ] <= 8'h00;
memory2_reg[899 ] <= 8'h00;
memory2_reg[900 ] <= 8'h00;
memory2_reg[901 ] <= 8'h00;
memory2_reg[902 ] <= 8'h00;
memory2_reg[903 ] <= 8'h00;
memory2_reg[904 ] <= 8'h00;
memory2_reg[905 ] <= 8'h00;
memory2_reg[906 ] <= 8'h00;
memory2_reg[907 ] <= 8'h00;
memory2_reg[908 ] <= 8'h00;
memory2_reg[909 ] <= 8'h00;
memory2_reg[910 ] <= 8'h00;
memory2_reg[911 ] <= 8'h00;
memory2_reg[912 ] <= 8'h00;
memory2_reg[913 ] <= 8'h00;
memory2_reg[914 ] <= 8'h00;
memory2_reg[915 ] <= 8'h00;
memory2_reg[916 ] <= 8'h00;
memory2_reg[917 ] <= 8'h00;
memory2_reg[918 ] <= 8'h00;
memory2_reg[919 ] <= 8'h00;
memory2_reg[920 ] <= 8'h00;
memory2_reg[921 ] <= 8'h00;
memory2_reg[922 ] <= 8'h00;
memory2_reg[923 ] <= 8'h00;
memory2_reg[924 ] <= 8'h00;
memory2_reg[925 ] <= 8'h00;
memory2_reg[926 ] <= 8'h00;
memory2_reg[927 ] <= 8'h00;
memory2_reg[928 ] <= 8'h00;
memory2_reg[929 ] <= 8'h00;
memory2_reg[930 ] <= 8'h00;
memory2_reg[931 ] <= 8'h00;
memory2_reg[932 ] <= 8'h00;
memory2_reg[933 ] <= 8'h00;
memory2_reg[934 ] <= 8'h00;
memory2_reg[935 ] <= 8'h00;
memory2_reg[936 ] <= 8'h00;
memory2_reg[937 ] <= 8'h00;
memory2_reg[938 ] <= 8'h00;
memory2_reg[939 ] <= 8'h00;
memory2_reg[940 ] <= 8'h00;
memory2_reg[941 ] <= 8'h00;
memory2_reg[942 ] <= 8'h00;
memory2_reg[943 ] <= 8'h00;
memory2_reg[944 ] <= 8'h00;
memory2_reg[945 ] <= 8'h00;
memory2_reg[946 ] <= 8'h00;
memory2_reg[947 ] <= 8'h00;
memory2_reg[948 ] <= 8'h00;
memory2_reg[949 ] <= 8'h00;
memory2_reg[950 ] <= 8'h00;
memory2_reg[951 ] <= 8'h00;
memory2_reg[952 ] <= 8'h00;
memory2_reg[953 ] <= 8'h00;
memory2_reg[954 ] <= 8'h00;
memory2_reg[955 ] <= 8'h00;
memory2_reg[956 ] <= 8'h00;
memory2_reg[957 ] <= 8'h00;
memory2_reg[958 ] <= 8'h00;
memory2_reg[959 ] <= 8'h00;
memory2_reg[960 ] <= 8'h00;
memory2_reg[961 ] <= 8'h00;
memory2_reg[962 ] <= 8'h00;
memory2_reg[963 ] <= 8'h00;
memory2_reg[964 ] <= 8'h00;
memory2_reg[965 ] <= 8'h00;
memory2_reg[966 ] <= 8'h00;
memory2_reg[967 ] <= 8'h00;
memory2_reg[968 ] <= 8'h00;
memory2_reg[969 ] <= 8'h00;
memory2_reg[970 ] <= 8'h00;
memory2_reg[971 ] <= 8'h00;
memory2_reg[972 ] <= 8'h00;
memory2_reg[973 ] <= 8'h00;
memory2_reg[974 ] <= 8'h00;
memory2_reg[975 ] <= 8'h00;
memory2_reg[976 ] <= 8'h00;
memory2_reg[977 ] <= 8'h00;
memory2_reg[978 ] <= 8'h00;
memory2_reg[979 ] <= 8'h00;
memory2_reg[980 ] <= 8'h00;
memory2_reg[981 ] <= 8'h00;
memory2_reg[982 ] <= 8'h00;
memory2_reg[983 ] <= 8'h00;
memory2_reg[984 ] <= 8'h00;
memory2_reg[985 ] <= 8'h00;
memory2_reg[986 ] <= 8'h00;
memory2_reg[987 ] <= 8'h00;
memory2_reg[988 ] <= 8'h00;
memory2_reg[989 ] <= 8'h00;
memory2_reg[990 ] <= 8'h00;
memory2_reg[991 ] <= 8'h00;
memory2_reg[992 ] <= 8'h00;
memory2_reg[993 ] <= 8'h00;
memory2_reg[994 ] <= 8'h00;
memory2_reg[995 ] <= 8'h00;
memory2_reg[996 ] <= 8'h00;
memory2_reg[997 ] <= 8'h00;
memory2_reg[998 ] <= 8'h00;
memory2_reg[999 ] <= 8'h00;
memory2_reg[1000] <= 8'h00;
memory2_reg[1001] <= 8'h00;
memory2_reg[1002] <= 8'h00;
memory2_reg[1003] <= 8'h00;
memory2_reg[1004] <= 8'h00;
memory2_reg[1005] <= 8'h00;
memory2_reg[1006] <= 8'h00;
memory2_reg[1007] <= 8'h00;
memory2_reg[1008] <= 8'h00;
memory2_reg[1009] <= 8'h00;
memory2_reg[1010] <= 8'h00;
memory2_reg[1011] <= 8'h00;
memory2_reg[1012] <= 8'h00;
memory2_reg[1013] <= 8'h00;
memory2_reg[1014] <= 8'h00;
memory2_reg[1015] <= 8'h00;
memory2_reg[1016] <= 8'h00;
memory2_reg[1017] <= 8'h00;
memory2_reg[1018] <= 8'h00;
memory2_reg[1019] <= 8'h00;
memory2_reg[1020] <= 8'h00;
memory2_reg[1021] <= 8'h00;
memory2_reg[1022] <= 8'h00;
memory2_reg[1023] <= 8'h00;

// Memory 3

memory3_reg[0   ] <= 8'h01;
memory3_reg[1   ] <= 8'h0F;
memory3_reg[2   ] <= 8'h02;
memory3_reg[3   ] <= 8'h0F;
memory3_reg[4   ] <= 8'h02;
memory3_reg[5   ] <= 8'h01;
memory3_reg[6   ] <= 8'h04;
memory3_reg[7   ] <= 8'h0F;
memory3_reg[8   ] <= 8'h05;
memory3_reg[9   ] <= 8'h01;
memory3_reg[10  ] <= 8'h01;
memory3_reg[11  ] <= 8'h0F;
memory3_reg[12  ] <= 8'h01;
memory3_reg[13  ] <= 8'h02;
memory3_reg[14  ] <= 8'h02;
memory3_reg[15  ] <= 8'h04;
memory3_reg[16  ] <= 8'h05;
memory3_reg[17  ] <= 8'h02;
memory3_reg[18  ] <= 8'h01;
memory3_reg[19  ] <= 8'h0F;
memory3_reg[20  ] <= 8'h02;
memory3_reg[21  ] <= 8'h0F;
memory3_reg[22  ] <= 8'h02;
memory3_reg[23  ] <= 8'h01;
memory3_reg[24  ] <= 8'h04;
memory3_reg[25  ] <= 8'h0F;
memory3_reg[26  ] <= 8'h05;
memory3_reg[27  ] <= 8'h01;
memory3_reg[28  ] <= 8'h01;
memory3_reg[29  ] <= 8'h0F;
memory3_reg[30  ] <= 8'h01;
memory3_reg[31  ] <= 8'h02;
memory3_reg[32  ] <= 8'h02;
memory3_reg[33  ] <= 8'h04;
memory3_reg[34  ] <= 8'h05;
memory3_reg[35  ] <= 8'h02;
memory3_reg[36  ] <= 8'h01;
memory3_reg[37  ] <= 8'h0F;
memory3_reg[38  ] <= 8'h02;
memory3_reg[39  ] <= 8'h0F;
memory3_reg[40  ] <= 8'h02;
memory3_reg[41  ] <= 8'h01;
memory3_reg[42  ] <= 8'h04;
memory3_reg[43  ] <= 8'h0F;
memory3_reg[44  ] <= 8'h05;
memory3_reg[45  ] <= 8'h01;
memory3_reg[46  ] <= 8'h01;
memory3_reg[47  ] <= 8'h0F;
memory3_reg[48  ] <= 8'h01;
memory3_reg[49  ] <= 8'h02;
memory3_reg[50  ] <= 8'h02;
memory3_reg[51  ] <= 8'h04;
memory3_reg[52  ] <= 8'h05;
memory3_reg[53  ] <= 8'h02;
memory3_reg[54  ] <= 8'h00;
memory3_reg[55  ] <= 8'h00;
memory3_reg[56  ] <= 8'h02;
memory3_reg[57  ] <= 8'h0F;
memory3_reg[58  ] <= 8'h02;
memory3_reg[59  ] <= 8'h0F;
memory3_reg[60  ] <= 8'h00;
memory3_reg[61  ] <= 8'h01;
memory3_reg[62  ] <= 8'h04;
memory3_reg[63  ] <= 8'h0F;
memory3_reg[64  ] <= 8'h05;
memory3_reg[65  ] <= 8'h02;
memory3_reg[66  ] <= 8'h02;
memory3_reg[67  ] <= 8'h0F;
memory3_reg[68  ] <= 8'h01;
memory3_reg[69  ] <= 8'h00;
memory3_reg[70  ] <= 8'h02;
memory3_reg[71  ] <= 8'h04;
memory3_reg[72  ] <= 8'h05;
memory3_reg[73  ] <= 8'h00;
memory3_reg[74  ] <= 8'h02;
memory3_reg[75  ] <= 8'h0F;
memory3_reg[76  ] <= 8'h02;
memory3_reg[77  ] <= 8'h0F;
memory3_reg[78  ] <= 8'h00;
memory3_reg[79  ] <= 8'h01;
memory3_reg[80  ] <= 8'h04;
memory3_reg[81  ] <= 8'h0F;
memory3_reg[82  ] <= 8'h05;
memory3_reg[83  ] <= 8'h02;
memory3_reg[84  ] <= 8'h02;
memory3_reg[85  ] <= 8'h0F;
memory3_reg[86  ] <= 8'h01;
memory3_reg[87  ] <= 8'h00;
memory3_reg[88  ] <= 8'h02;
memory3_reg[89  ] <= 8'h04;
memory3_reg[90  ] <= 8'h05;
memory3_reg[91  ] <= 8'h00;
memory3_reg[92  ] <= 8'h02;
memory3_reg[93  ] <= 8'h0F;
memory3_reg[94  ] <= 8'h02;
memory3_reg[95  ] <= 8'h0F;
memory3_reg[96  ] <= 8'h00;
memory3_reg[97  ] <= 8'h01;
memory3_reg[98  ] <= 8'h04;
memory3_reg[99  ] <= 8'h0F;
memory3_reg[100 ] <= 8'h05;
memory3_reg[101 ] <= 8'h02;
memory3_reg[102 ] <= 8'h02;
memory3_reg[103 ] <= 8'h0F;
memory3_reg[104 ] <= 8'h01;
memory3_reg[105 ] <= 8'h00;
memory3_reg[106 ] <= 8'h02;
memory3_reg[107 ] <= 8'h04;
memory3_reg[108 ] <= 8'h05;
memory3_reg[109 ] <= 8'h00;
memory3_reg[110 ] <= 8'h00;
memory3_reg[111 ] <= 8'h00;
memory3_reg[112 ] <= 8'h00;
memory3_reg[113 ] <= 8'h0F;
memory3_reg[114 ] <= 8'h02;
memory3_reg[115 ] <= 8'h0F;
memory3_reg[116 ] <= 8'h01;
memory3_reg[117 ] <= 8'h01;
memory3_reg[118 ] <= 8'h04;
memory3_reg[119 ] <= 8'h0F;
memory3_reg[120 ] <= 8'h05;
memory3_reg[121 ] <= 8'h00;
memory3_reg[122 ] <= 8'h00;
memory3_reg[123 ] <= 8'h0F;
memory3_reg[124 ] <= 8'h01;
memory3_reg[125 ] <= 8'h01;
memory3_reg[126 ] <= 8'h02;
memory3_reg[127 ] <= 8'h04;
memory3_reg[128 ] <= 8'h05;
memory3_reg[129 ] <= 8'h01;
memory3_reg[130 ] <= 8'h00;
memory3_reg[131 ] <= 8'h0F;
memory3_reg[132 ] <= 8'h02;
memory3_reg[133 ] <= 8'h0F;
memory3_reg[134 ] <= 8'h01;
memory3_reg[135 ] <= 8'h01;
memory3_reg[136 ] <= 8'h04;
memory3_reg[137 ] <= 8'h0F;
memory3_reg[138 ] <= 8'h05;
memory3_reg[139 ] <= 8'h00;
memory3_reg[140 ] <= 8'h00;
memory3_reg[141 ] <= 8'h0F;
memory3_reg[142 ] <= 8'h01;
memory3_reg[143 ] <= 8'h01;
memory3_reg[144 ] <= 8'h02;
memory3_reg[145 ] <= 8'h04;
memory3_reg[146 ] <= 8'h05;
memory3_reg[147 ] <= 8'h01;
memory3_reg[148 ] <= 8'h00;
memory3_reg[149 ] <= 8'h0F;
memory3_reg[150 ] <= 8'h02;
memory3_reg[151 ] <= 8'h0F;
memory3_reg[152 ] <= 8'h01;
memory3_reg[153 ] <= 8'h01;
memory3_reg[154 ] <= 8'h04;
memory3_reg[155 ] <= 8'h0F;
memory3_reg[156 ] <= 8'h05;
memory3_reg[157 ] <= 8'h00;
memory3_reg[158 ] <= 8'h00;
memory3_reg[159 ] <= 8'h0F;
memory3_reg[160 ] <= 8'h01;
memory3_reg[161 ] <= 8'h01;
memory3_reg[162 ] <= 8'h02;
memory3_reg[163 ] <= 8'h04;
memory3_reg[164 ] <= 8'h05;
memory3_reg[165 ] <= 8'h01;
memory3_reg[166 ] <= 8'h00;
memory3_reg[167 ] <= 8'h00;
memory3_reg[168 ] <= 8'h00;
memory3_reg[169 ] <= 8'h00;
memory3_reg[170 ] <= 8'h04;
memory3_reg[171 ] <= 8'h01;
memory3_reg[172 ] <= 8'h01;
memory3_reg[173 ] <= 8'h08;
memory3_reg[174 ] <= 8'h02;
memory3_reg[175 ] <= 8'h02;
memory3_reg[176 ] <= 8'h0C;
memory3_reg[177 ] <= 8'h00;
memory3_reg[178 ] <= 8'h00;
memory3_reg[179 ] <= 8'h00;
memory3_reg[180 ] <= 8'h05;
memory3_reg[181 ] <= 8'h01;
memory3_reg[182 ] <= 8'h01;
memory3_reg[183 ] <= 8'h09;
memory3_reg[184 ] <= 8'h02;
memory3_reg[185 ] <= 8'h02;
memory3_reg[186 ] <= 8'h0D;
memory3_reg[187 ] <= 8'h01;
memory3_reg[188 ] <= 8'h00;
memory3_reg[189 ] <= 8'h00;
memory3_reg[190 ] <= 8'h06;
memory3_reg[191 ] <= 8'h01;
memory3_reg[192 ] <= 8'h01;
memory3_reg[193 ] <= 8'h0A;
memory3_reg[194 ] <= 8'h02;
memory3_reg[195 ] <= 8'h02;
memory3_reg[196 ] <= 8'h0E;
memory3_reg[197 ] <= 8'h02;
memory3_reg[198 ] <= 8'h00;
memory3_reg[199 ] <= 8'h00;
memory3_reg[200 ] <= 8'h00;
memory3_reg[201 ] <= 8'h00;
memory3_reg[202 ] <= 8'h00;
memory3_reg[203 ] <= 8'h00;
memory3_reg[204 ] <= 8'h00;
memory3_reg[205 ] <= 8'h00;
memory3_reg[206 ] <= 8'h00;
memory3_reg[207 ] <= 8'h00;
memory3_reg[208 ] <= 8'h00;
memory3_reg[209 ] <= 8'h00;
memory3_reg[210 ] <= 8'h00;
memory3_reg[211 ] <= 8'h00;
memory3_reg[212 ] <= 8'h00;
memory3_reg[213 ] <= 8'h00;
memory3_reg[214 ] <= 8'h00;
memory3_reg[215 ] <= 8'h00;
memory3_reg[216 ] <= 8'h00;
memory3_reg[217 ] <= 8'h00;
memory3_reg[218 ] <= 8'h00;
memory3_reg[219 ] <= 8'h00;
memory3_reg[220 ] <= 8'h00;
memory3_reg[221 ] <= 8'h00;
memory3_reg[222 ] <= 8'h00;
memory3_reg[223 ] <= 8'h00;
memory3_reg[224 ] <= 8'h00;
memory3_reg[225 ] <= 8'h00;
memory3_reg[226 ] <= 8'h00;
memory3_reg[227 ] <= 8'h00;
memory3_reg[228 ] <= 8'h00;
memory3_reg[229 ] <= 8'h00;
memory3_reg[230 ] <= 8'h00;
memory3_reg[231 ] <= 8'h00;
memory3_reg[232 ] <= 8'h00;
memory3_reg[233 ] <= 8'h00;
memory3_reg[234 ] <= 8'h00;
memory3_reg[235 ] <= 8'h00;
memory3_reg[236 ] <= 8'h00;
memory3_reg[237 ] <= 8'h00;
memory3_reg[238 ] <= 8'h00;
memory3_reg[239 ] <= 8'h00;
memory3_reg[240 ] <= 8'h00;
memory3_reg[241 ] <= 8'h00;
memory3_reg[242 ] <= 8'h00;
memory3_reg[243 ] <= 8'h00;
memory3_reg[244 ] <= 8'h00;
memory3_reg[245 ] <= 8'h00;
memory3_reg[246 ] <= 8'h00;
memory3_reg[247 ] <= 8'h00;
memory3_reg[248 ] <= 8'h00;
memory3_reg[249 ] <= 8'h00;
memory3_reg[250 ] <= 8'h00;
memory3_reg[251 ] <= 8'h00;
memory3_reg[252 ] <= 8'h00;
memory3_reg[253 ] <= 8'h00;
memory3_reg[254 ] <= 8'h00;
memory3_reg[255 ] <= 8'h00;
memory3_reg[256 ] <= 8'h0F;
memory3_reg[257 ] <= 8'h04;
memory3_reg[258 ] <= 8'h04;
memory3_reg[259 ] <= 8'h08;
memory3_reg[260 ] <= 8'h08;
memory3_reg[261 ] <= 8'h0C;
memory3_reg[262 ] <= 8'h0C;
memory3_reg[263 ] <= 8'h03;
memory3_reg[264 ] <= 8'h04;
memory3_reg[265 ] <= 8'h05;
memory3_reg[266 ] <= 8'h08;
memory3_reg[267 ] <= 8'h09;
memory3_reg[268 ] <= 8'h0C;
memory3_reg[269 ] <= 8'h0D;
memory3_reg[270 ] <= 8'h04;
memory3_reg[271 ] <= 8'h04;
memory3_reg[272 ] <= 8'h06;
memory3_reg[273 ] <= 8'h08;
memory3_reg[274 ] <= 8'h0A;
memory3_reg[275 ] <= 8'h0C;
memory3_reg[276 ] <= 8'h0E;
memory3_reg[277 ] <= 8'h05;
memory3_reg[278 ] <= 8'h05;
memory3_reg[279 ] <= 8'h04;
memory3_reg[280 ] <= 8'h09;
memory3_reg[281 ] <= 8'h08;
memory3_reg[282 ] <= 8'h0D;
memory3_reg[283 ] <= 8'h0C;
memory3_reg[284 ] <= 8'h06;
memory3_reg[285 ] <= 8'h05;
memory3_reg[286 ] <= 8'h05;
memory3_reg[287 ] <= 8'h09;
memory3_reg[288 ] <= 8'h09;
memory3_reg[289 ] <= 8'h0D;
memory3_reg[290 ] <= 8'h0D;
memory3_reg[291 ] <= 8'h07;
memory3_reg[292 ] <= 8'h05;
memory3_reg[293 ] <= 8'h06;
memory3_reg[294 ] <= 8'h09;
memory3_reg[295 ] <= 8'h0A;
memory3_reg[296 ] <= 8'h0D;
memory3_reg[297 ] <= 8'h0E;
memory3_reg[298 ] <= 8'h08;
memory3_reg[299 ] <= 8'h06;
memory3_reg[300 ] <= 8'h04;
memory3_reg[301 ] <= 8'h0A;
memory3_reg[302 ] <= 8'h08;
memory3_reg[303 ] <= 8'h0E;
memory3_reg[304 ] <= 8'h0C;
memory3_reg[305 ] <= 8'h09;
memory3_reg[306 ] <= 8'h06;
memory3_reg[307 ] <= 8'h05;
memory3_reg[308 ] <= 8'h0A;
memory3_reg[309 ] <= 8'h09;
memory3_reg[310 ] <= 8'h0E;
memory3_reg[311 ] <= 8'h0D;
memory3_reg[312 ] <= 8'h0A;
memory3_reg[313 ] <= 8'h06;
memory3_reg[314 ] <= 8'h06;
memory3_reg[315 ] <= 8'h0A;
memory3_reg[316 ] <= 8'h0A;
memory3_reg[317 ] <= 8'h0E;
memory3_reg[318 ] <= 8'h0E;
memory3_reg[319 ] <= 8'h0B;
memory3_reg[320 ] <= 8'h0F;
memory3_reg[321 ] <= 8'h0C;
memory3_reg[322 ] <= 8'h00;
memory3_reg[323 ] <= 8'h03;
memory3_reg[324 ] <= 8'h01;
memory3_reg[325 ] <= 8'h06;
memory3_reg[326 ] <= 8'h02;
memory3_reg[327 ] <= 8'h09;
memory3_reg[328 ] <= 8'h00;
memory3_reg[329 ] <= 8'h0D;
memory3_reg[330 ] <= 8'h00;
memory3_reg[331 ] <= 8'h04;
memory3_reg[332 ] <= 8'h01;
memory3_reg[333 ] <= 8'h07;
memory3_reg[334 ] <= 8'h02;
memory3_reg[335 ] <= 8'h0A;
memory3_reg[336 ] <= 8'h01;
memory3_reg[337 ] <= 8'h0E;
memory3_reg[338 ] <= 8'h00;
memory3_reg[339 ] <= 8'h05;
memory3_reg[340 ] <= 8'h01;
memory3_reg[341 ] <= 8'h08;
memory3_reg[342 ] <= 8'h02;
memory3_reg[343 ] <= 8'h0B;
memory3_reg[344 ] <= 8'h02;
memory3_reg[345 ] <= 8'h00;
memory3_reg[346 ] <= 8'h06;
memory3_reg[347 ] <= 8'h07;
memory3_reg[348 ] <= 8'h0F;
memory3_reg[349 ] <= 8'h00;
memory3_reg[350 ] <= 8'h00;
memory3_reg[351 ] <= 8'h00;
memory3_reg[352 ] <= 8'h0F;
memory3_reg[353 ] <= 8'h00;
memory3_reg[354 ] <= 8'h00;
memory3_reg[355 ] <= 8'h00;
memory3_reg[356 ] <= 8'h0F;
memory3_reg[357 ] <= 8'h00;
memory3_reg[358 ] <= 8'h00;
memory3_reg[359 ] <= 8'h00;
memory3_reg[360 ] <= 8'h00;
memory3_reg[361 ] <= 8'h00;
memory3_reg[362 ] <= 8'h00;
memory3_reg[363 ] <= 8'h00;
memory3_reg[364 ] <= 8'h00;
memory3_reg[365 ] <= 8'h00;
memory3_reg[366 ] <= 8'h00;
memory3_reg[367 ] <= 8'h00;
memory3_reg[368 ] <= 8'h00;
memory3_reg[369 ] <= 8'h01;
memory3_reg[370 ] <= 8'h00;
memory3_reg[371 ] <= 8'h00;
memory3_reg[372 ] <= 8'h0C;
memory3_reg[373 ] <= 8'h0D;
memory3_reg[374 ] <= 8'h0E;
memory3_reg[375 ] <= 8'h00;
memory3_reg[376 ] <= 8'h0C;
memory3_reg[377 ] <= 8'h0D;
memory3_reg[378 ] <= 8'h0E;
memory3_reg[379 ] <= 8'h00;
memory3_reg[380 ] <= 8'h00;
memory3_reg[381 ] <= 8'h0F;
memory3_reg[382 ] <= 8'h00;
memory3_reg[383 ] <= 8'h00;
memory3_reg[384 ] <= 8'h0F;
memory3_reg[385 ] <= 8'h00;
memory3_reg[386 ] <= 8'h00;
memory3_reg[387 ] <= 8'h04;
memory3_reg[388 ] <= 8'h01;
memory3_reg[389 ] <= 8'h05;
memory3_reg[390 ] <= 8'h02;
memory3_reg[391 ] <= 8'h06;
memory3_reg[392 ] <= 8'h00;
memory3_reg[393 ] <= 8'h01;
memory3_reg[394 ] <= 8'h00;
memory3_reg[395 ] <= 8'h08;
memory3_reg[396 ] <= 8'h01;
memory3_reg[397 ] <= 8'h09;
memory3_reg[398 ] <= 8'h02;
memory3_reg[399 ] <= 8'h0A;
memory3_reg[400 ] <= 8'h01;
memory3_reg[401 ] <= 8'h02;
memory3_reg[402 ] <= 8'h00;
memory3_reg[403 ] <= 8'h0C;
memory3_reg[404 ] <= 8'h01;
memory3_reg[405 ] <= 8'h0D;
memory3_reg[406 ] <= 8'h02;
memory3_reg[407 ] <= 8'h0E;
memory3_reg[408 ] <= 8'h02;
memory3_reg[409 ] <= 8'h00;
memory3_reg[410 ] <= 8'h00;
memory3_reg[411 ] <= 8'h00;
memory3_reg[412 ] <= 8'h00;
memory3_reg[413 ] <= 8'h00;
memory3_reg[414 ] <= 8'h00;
memory3_reg[415 ] <= 8'h0C;
memory3_reg[416 ] <= 8'h0C;
memory3_reg[417 ] <= 8'h0F;
memory3_reg[418 ] <= 8'h03;
memory3_reg[419 ] <= 8'h0C;
memory3_reg[420 ] <= 8'h01;
memory3_reg[421 ] <= 8'h01;
memory3_reg[422 ] <= 8'h00;
memory3_reg[423 ] <= 8'h0D;
memory3_reg[424 ] <= 8'h0D;
memory3_reg[425 ] <= 8'h0F;
memory3_reg[426 ] <= 8'h03;
memory3_reg[427 ] <= 8'h0D;
memory3_reg[428 ] <= 8'h02;
memory3_reg[429 ] <= 8'h02;
memory3_reg[430 ] <= 8'h00;
memory3_reg[431 ] <= 8'h0E;
memory3_reg[432 ] <= 8'h0E;
memory3_reg[433 ] <= 8'h0F;
memory3_reg[434 ] <= 8'h03;
memory3_reg[435 ] <= 8'h0E;
memory3_reg[436 ] <= 8'h0F;
memory3_reg[437 ] <= 8'h0C;
memory3_reg[438 ] <= 8'h04;
memory3_reg[439 ] <= 8'h0D;
memory3_reg[440 ] <= 8'h08;
memory3_reg[441 ] <= 8'h0E;
memory3_reg[442 ] <= 8'h0C;
memory3_reg[443 ] <= 8'h00;
memory3_reg[444 ] <= 8'h0C;
memory3_reg[445 ] <= 8'h05;
memory3_reg[446 ] <= 8'h0D;
memory3_reg[447 ] <= 8'h09;
memory3_reg[448 ] <= 8'h0E;
memory3_reg[449 ] <= 8'h0D;
memory3_reg[450 ] <= 8'h01;
memory3_reg[451 ] <= 8'h0C;
memory3_reg[452 ] <= 8'h06;
memory3_reg[453 ] <= 8'h0D;
memory3_reg[454 ] <= 8'h0A;
memory3_reg[455 ] <= 8'h0E;
memory3_reg[456 ] <= 8'h0E;
memory3_reg[457 ] <= 8'h02;
memory3_reg[458 ] <= 8'h00;
memory3_reg[459 ] <= 8'h06;
memory3_reg[460 ] <= 8'h07;
memory3_reg[461 ] <= 8'h07;
memory3_reg[462 ] <= 8'h07;
memory3_reg[463 ] <= 8'h0B;
memory3_reg[464 ] <= 8'h00;
memory3_reg[465 ] <= 8'h00;
memory3_reg[466 ] <= 8'h08;
memory3_reg[467 ] <= 8'h01;
memory3_reg[468 ] <= 8'h01;
memory3_reg[469 ] <= 8'h09;
memory3_reg[470 ] <= 8'h02;
memory3_reg[471 ] <= 8'h02;
memory3_reg[472 ] <= 8'h0A;
memory3_reg[473 ] <= 8'h00;
memory3_reg[474 ] <= 8'h00;
memory3_reg[475 ] <= 8'h00;
memory3_reg[476 ] <= 8'h00;
memory3_reg[477 ] <= 8'h04;
memory3_reg[478 ] <= 8'h01;
memory3_reg[479 ] <= 8'h05;
memory3_reg[480 ] <= 8'h02;
memory3_reg[481 ] <= 8'h06;
memory3_reg[482 ] <= 8'h00;
memory3_reg[483 ] <= 8'h08;
memory3_reg[484 ] <= 8'h01;
memory3_reg[485 ] <= 8'h09;
memory3_reg[486 ] <= 8'h02;
memory3_reg[487 ] <= 8'h0A;
memory3_reg[488 ] <= 8'h00;
memory3_reg[489 ] <= 8'h0C;
memory3_reg[490 ] <= 8'h01;
memory3_reg[491 ] <= 8'h0D;
memory3_reg[492 ] <= 8'h02;
memory3_reg[493 ] <= 8'h0E;
memory3_reg[494 ] <= 8'h00;
memory3_reg[495 ] <= 8'h00;
memory3_reg[496 ] <= 8'h01;
memory3_reg[497 ] <= 8'h01;
memory3_reg[498 ] <= 8'h02;
memory3_reg[499 ] <= 8'h02;
memory3_reg[500 ] <= 8'h00;
memory3_reg[501 ] <= 8'h00;
memory3_reg[502 ] <= 8'h00;
memory3_reg[503 ] <= 8'h00;
memory3_reg[504 ] <= 8'h00;
memory3_reg[505 ] <= 8'h00;
memory3_reg[506 ] <= 8'h00;
memory3_reg[507 ] <= 8'h00;
memory3_reg[508 ] <= 8'h00;
memory3_reg[509 ] <= 8'h00;
memory3_reg[510 ] <= 8'h00;
memory3_reg[511 ] <= 8'h00;
memory3_reg[512 ] <= 8'h00;
memory3_reg[513 ] <= 8'h04;
memory3_reg[514 ] <= 8'h01;
memory3_reg[515 ] <= 8'h05;
memory3_reg[516 ] <= 8'h02;
memory3_reg[517 ] <= 8'h06;
memory3_reg[518 ] <= 8'h00;
memory3_reg[519 ] <= 8'h08;
memory3_reg[520 ] <= 8'h01;
memory3_reg[521 ] <= 8'h09;
memory3_reg[522 ] <= 8'h02;
memory3_reg[523 ] <= 8'h0A;
memory3_reg[524 ] <= 8'h00;
memory3_reg[525 ] <= 8'h0C;
memory3_reg[526 ] <= 8'h01;
memory3_reg[527 ] <= 8'h0D;
memory3_reg[528 ] <= 8'h02;
memory3_reg[529 ] <= 8'h0E;
memory3_reg[530 ] <= 8'h00;
memory3_reg[531 ] <= 8'h00;
memory3_reg[532 ] <= 8'h01;
memory3_reg[533 ] <= 8'h01;
memory3_reg[534 ] <= 8'h02;
memory3_reg[535 ] <= 8'h02;
memory3_reg[536 ] <= 8'h0F;
memory3_reg[537 ] <= 8'h01;
memory3_reg[538 ] <= 8'h00;
memory3_reg[539 ] <= 8'h01;
memory3_reg[540 ] <= 8'h02;
memory3_reg[541 ] <= 8'h00;
memory3_reg[542 ] <= 8'h02;
memory3_reg[543 ] <= 8'h00;
memory3_reg[544 ] <= 8'h0F;
memory3_reg[545 ] <= 8'h04;
memory3_reg[546 ] <= 8'h04;
memory3_reg[547 ] <= 8'h08;
memory3_reg[548 ] <= 8'h08;
memory3_reg[549 ] <= 8'h0C;
memory3_reg[550 ] <= 8'h00;
memory3_reg[551 ] <= 8'h00;
memory3_reg[552 ] <= 8'h0C;
memory3_reg[553 ] <= 8'h0D;
memory3_reg[554 ] <= 8'h0D;
memory3_reg[555 ] <= 8'h0D;
memory3_reg[556 ] <= 8'h08;
memory3_reg[557 ] <= 8'h0F;
memory3_reg[558 ] <= 8'h0D;
memory3_reg[559 ] <= 8'h04;
memory3_reg[560 ] <= 8'h0E;
memory3_reg[561 ] <= 8'h04;
memory3_reg[562 ] <= 8'h0F;
memory3_reg[563 ] <= 8'h06;
memory3_reg[564 ] <= 8'h0F;
memory3_reg[565 ] <= 8'h08;
memory3_reg[566 ] <= 8'h0A;
memory3_reg[567 ] <= 8'h0E;
memory3_reg[568 ] <= 8'h0A;
memory3_reg[569 ] <= 8'h08;
memory3_reg[570 ] <= 8'h04;
memory3_reg[571 ] <= 8'h0F;
memory3_reg[572 ] <= 8'h05;
memory3_reg[573 ] <= 8'h0F;
memory3_reg[574 ] <= 8'h08;
memory3_reg[575 ] <= 8'h09;
memory3_reg[576 ] <= 8'h0E;
memory3_reg[577 ] <= 8'h09;
memory3_reg[578 ] <= 8'h09;
memory3_reg[579 ] <= 8'h04;
memory3_reg[580 ] <= 8'h06;
memory3_reg[581 ] <= 8'h0F;
memory3_reg[582 ] <= 8'h06;
memory3_reg[583 ] <= 8'h08;
memory3_reg[584 ] <= 8'h0E;
memory3_reg[585 ] <= 8'h0A;
memory3_reg[586 ] <= 8'h0A;
memory3_reg[587 ] <= 8'h0F;
memory3_reg[588 ] <= 8'h04;
memory3_reg[589 ] <= 8'h05;
memory3_reg[590 ] <= 8'h0F;
memory3_reg[591 ] <= 8'h05;
memory3_reg[592 ] <= 8'h08;
memory3_reg[593 ] <= 8'h0E;
memory3_reg[594 ] <= 8'h09;
memory3_reg[595 ] <= 8'h0B;
memory3_reg[596 ] <= 8'h0F;
memory3_reg[597 ] <= 8'h0F;
memory3_reg[598 ] <= 8'h01;
memory3_reg[599 ] <= 8'h0F;
memory3_reg[600 ] <= 8'h0F;
memory3_reg[601 ] <= 8'h07;
memory3_reg[602 ] <= 8'h06;
memory3_reg[603 ] <= 8'h0B;
memory3_reg[604 ] <= 8'h0A;
memory3_reg[605 ] <= 8'h0F;
memory3_reg[606 ] <= 8'h0E;
memory3_reg[607 ] <= 8'h0C;
memory3_reg[608 ] <= 8'h0F;
memory3_reg[609 ] <= 8'h04;
memory3_reg[610 ] <= 8'h00;
memory3_reg[611 ] <= 8'h07;
memory3_reg[612 ] <= 8'h0C;
memory3_reg[613 ] <= 8'h06;
memory3_reg[614 ] <= 8'h03;
memory3_reg[615 ] <= 8'h0F;
memory3_reg[616 ] <= 8'h08;
memory3_reg[617 ] <= 8'h00;
memory3_reg[618 ] <= 8'h0B;
memory3_reg[619 ] <= 8'h0C;
memory3_reg[620 ] <= 8'h0A;
memory3_reg[621 ] <= 8'h07;
memory3_reg[622 ] <= 8'h03;
memory3_reg[623 ] <= 8'h0F;
memory3_reg[624 ] <= 8'h0C;
memory3_reg[625 ] <= 8'h00;
memory3_reg[626 ] <= 8'h0F;
memory3_reg[627 ] <= 8'h0C;
memory3_reg[628 ] <= 8'h0E;
memory3_reg[629 ] <= 8'h0B;
memory3_reg[630 ] <= 8'h00;
memory3_reg[631 ] <= 8'h00;
memory3_reg[632 ] <= 8'h0F;
memory3_reg[633 ] <= 8'h0F;
memory3_reg[634 ] <= 8'h01;
memory3_reg[635 ] <= 8'h0F;
memory3_reg[636 ] <= 8'h0F;
memory3_reg[637 ] <= 8'h06;
memory3_reg[638 ] <= 8'h00;
memory3_reg[639 ] <= 8'h07;
memory3_reg[640 ] <= 8'h03;
memory3_reg[641 ] <= 8'h0F;
memory3_reg[642 ] <= 8'h0A;
memory3_reg[643 ] <= 8'h00;
memory3_reg[644 ] <= 8'h0B;
memory3_reg[645 ] <= 8'h07;
memory3_reg[646 ] <= 8'h03;
memory3_reg[647 ] <= 8'h0F;
memory3_reg[648 ] <= 8'h0E;
memory3_reg[649 ] <= 8'h00;
memory3_reg[650 ] <= 8'h0F;
memory3_reg[651 ] <= 8'h0B;
memory3_reg[652 ] <= 8'h0F;
memory3_reg[653 ] <= 8'h0F;
memory3_reg[654 ] <= 8'h01;
memory3_reg[655 ] <= 8'h0F;
memory3_reg[656 ] <= 8'h0F;
memory3_reg[657 ] <= 8'h07;
memory3_reg[658 ] <= 8'h06;
memory3_reg[659 ] <= 8'h0B;
memory3_reg[660 ] <= 8'h0A;
memory3_reg[661 ] <= 8'h0F;
memory3_reg[662 ] <= 8'h0E;
memory3_reg[663 ] <= 8'h0C;
memory3_reg[664 ] <= 8'h0F;
memory3_reg[665 ] <= 8'h0F;
memory3_reg[666 ] <= 8'h06;
memory3_reg[667 ] <= 8'h00;
memory3_reg[668 ] <= 8'h07;
memory3_reg[669 ] <= 8'h0C;
memory3_reg[670 ] <= 8'h06;
memory3_reg[671 ] <= 8'h03;
memory3_reg[672 ] <= 8'h0F;
memory3_reg[673 ] <= 8'h0A;
memory3_reg[674 ] <= 8'h00;
memory3_reg[675 ] <= 8'h0B;
memory3_reg[676 ] <= 8'h0C;
memory3_reg[677 ] <= 8'h0A;
memory3_reg[678 ] <= 8'h07;
memory3_reg[679 ] <= 8'h03;
memory3_reg[680 ] <= 8'h0F;
memory3_reg[681 ] <= 8'h0E;
memory3_reg[682 ] <= 8'h00;
memory3_reg[683 ] <= 8'h0F;
memory3_reg[684 ] <= 8'h0C;
memory3_reg[685 ] <= 8'h0E;
memory3_reg[686 ] <= 8'h0B;
memory3_reg[687 ] <= 8'h00;
memory3_reg[688 ] <= 8'h0F;
memory3_reg[689 ] <= 8'h07;
memory3_reg[690 ] <= 8'h04;
memory3_reg[691 ] <= 8'h0B;
memory3_reg[692 ] <= 8'h08;
memory3_reg[693 ] <= 8'h0F;
memory3_reg[694 ] <= 8'h0C;
memory3_reg[695 ] <= 8'h0F;
memory3_reg[696 ] <= 8'h00;
memory3_reg[697 ] <= 8'h01;
memory3_reg[698 ] <= 8'h0D;
memory3_reg[699 ] <= 8'h02;
memory3_reg[700 ] <= 8'h01;
memory3_reg[701 ] <= 8'h02;
memory3_reg[702 ] <= 8'h0D;
memory3_reg[703 ] <= 8'h03;
memory3_reg[704 ] <= 8'h03;
memory3_reg[705 ] <= 8'h00;
memory3_reg[706 ] <= 8'h00;
memory3_reg[707 ] <= 8'h0C;
memory3_reg[708 ] <= 8'h00;
memory3_reg[709 ] <= 8'h00;
memory3_reg[710 ] <= 8'h00;
memory3_reg[711 ] <= 8'h00;
memory3_reg[712 ] <= 8'h00;
memory3_reg[713 ] <= 8'h00;
memory3_reg[714 ] <= 8'h00;
memory3_reg[715 ] <= 8'h00;
memory3_reg[716 ] <= 8'h00;
memory3_reg[717 ] <= 8'h00;
memory3_reg[718 ] <= 8'h00;
memory3_reg[719 ] <= 8'h00;
memory3_reg[720 ] <= 8'h00;
memory3_reg[721 ] <= 8'h00;
memory3_reg[722 ] <= 8'h00;
memory3_reg[723 ] <= 8'h00;
memory3_reg[724 ] <= 8'h00;
memory3_reg[725 ] <= 8'h00;
memory3_reg[726 ] <= 8'h00;
memory3_reg[727 ] <= 8'h00;
memory3_reg[728 ] <= 8'h00;
memory3_reg[729 ] <= 8'h00;
memory3_reg[730 ] <= 8'h00;
memory3_reg[731 ] <= 8'h00;
memory3_reg[732 ] <= 8'h00;
memory3_reg[733 ] <= 8'h00;
memory3_reg[734 ] <= 8'h00;
memory3_reg[735 ] <= 8'h00;
memory3_reg[736 ] <= 8'h00;
memory3_reg[737 ] <= 8'h00;
memory3_reg[738 ] <= 8'h00;
memory3_reg[739 ] <= 8'h00;
memory3_reg[740 ] <= 8'h00;
memory3_reg[741 ] <= 8'h00;
memory3_reg[742 ] <= 8'h00;
memory3_reg[743 ] <= 8'h00;
memory3_reg[744 ] <= 8'h00;
memory3_reg[745 ] <= 8'h00;
memory3_reg[746 ] <= 8'h00;
memory3_reg[747 ] <= 8'h00;
memory3_reg[748 ] <= 8'h00;
memory3_reg[749 ] <= 8'h00;
memory3_reg[750 ] <= 8'h00;
memory3_reg[751 ] <= 8'h00;
memory3_reg[752 ] <= 8'h00;
memory3_reg[753 ] <= 8'h00;
memory3_reg[754 ] <= 8'h00;
memory3_reg[755 ] <= 8'h00;
memory3_reg[756 ] <= 8'h00;
memory3_reg[757 ] <= 8'h00;
memory3_reg[758 ] <= 8'h00;
memory3_reg[759 ] <= 8'h00;
memory3_reg[760 ] <= 8'h00;
memory3_reg[761 ] <= 8'h00;
memory3_reg[762 ] <= 8'h00;
memory3_reg[763 ] <= 8'h00;
memory3_reg[764 ] <= 8'h00;
memory3_reg[765 ] <= 8'h00;
memory3_reg[766 ] <= 8'h00;
memory3_reg[767 ] <= 8'h00;
memory3_reg[768 ] <= 8'h00;
memory3_reg[769 ] <= 8'h00;
memory3_reg[770 ] <= 8'h00;
memory3_reg[771 ] <= 8'h00;
memory3_reg[772 ] <= 8'h00;
memory3_reg[773 ] <= 8'h00;
memory3_reg[774 ] <= 8'h00;
memory3_reg[775 ] <= 8'h00;
memory3_reg[776 ] <= 8'h00;
memory3_reg[777 ] <= 8'h00;
memory3_reg[778 ] <= 8'h00;
memory3_reg[779 ] <= 8'h00;
memory3_reg[780 ] <= 8'h00;
memory3_reg[781 ] <= 8'h00;
memory3_reg[782 ] <= 8'h00;
memory3_reg[783 ] <= 8'h00;
memory3_reg[784 ] <= 8'h00;
memory3_reg[785 ] <= 8'h00;
memory3_reg[786 ] <= 8'h00;
memory3_reg[787 ] <= 8'h00;
memory3_reg[788 ] <= 8'h00;
memory3_reg[789 ] <= 8'h00;
memory3_reg[790 ] <= 8'h00;
memory3_reg[791 ] <= 8'h00;
memory3_reg[792 ] <= 8'h00;
memory3_reg[793 ] <= 8'h00;
memory3_reg[794 ] <= 8'h00;
memory3_reg[795 ] <= 8'h00;
memory3_reg[796 ] <= 8'h00;
memory3_reg[797 ] <= 8'h00;
memory3_reg[798 ] <= 8'h00;
memory3_reg[799 ] <= 8'h00;
memory3_reg[800 ] <= 8'h00;
memory3_reg[801 ] <= 8'h00;
memory3_reg[802 ] <= 8'h00;
memory3_reg[803 ] <= 8'h00;
memory3_reg[804 ] <= 8'h00;
memory3_reg[805 ] <= 8'h00;
memory3_reg[806 ] <= 8'h00;
memory3_reg[807 ] <= 8'h00;
memory3_reg[808 ] <= 8'h00;
memory3_reg[809 ] <= 8'h00;
memory3_reg[810 ] <= 8'h00;
memory3_reg[811 ] <= 8'h00;
memory3_reg[812 ] <= 8'h00;
memory3_reg[813 ] <= 8'h00;
memory3_reg[814 ] <= 8'h00;
memory3_reg[815 ] <= 8'h00;
memory3_reg[816 ] <= 8'h00;
memory3_reg[817 ] <= 8'h00;
memory3_reg[818 ] <= 8'h00;
memory3_reg[819 ] <= 8'h00;
memory3_reg[820 ] <= 8'h00;
memory3_reg[821 ] <= 8'h00;
memory3_reg[822 ] <= 8'h00;
memory3_reg[823 ] <= 8'h00;
memory3_reg[824 ] <= 8'h00;
memory3_reg[825 ] <= 8'h00;
memory3_reg[826 ] <= 8'h00;
memory3_reg[827 ] <= 8'h00;
memory3_reg[828 ] <= 8'h00;
memory3_reg[829 ] <= 8'h00;
memory3_reg[830 ] <= 8'h00;
memory3_reg[831 ] <= 8'h00;
memory3_reg[832 ] <= 8'h00;
memory3_reg[833 ] <= 8'h00;
memory3_reg[834 ] <= 8'h00;
memory3_reg[835 ] <= 8'h00;
memory3_reg[836 ] <= 8'h00;
memory3_reg[837 ] <= 8'h00;
memory3_reg[838 ] <= 8'h00;
memory3_reg[839 ] <= 8'h00;
memory3_reg[840 ] <= 8'h00;
memory3_reg[841 ] <= 8'h00;
memory3_reg[842 ] <= 8'h00;
memory3_reg[843 ] <= 8'h00;
memory3_reg[844 ] <= 8'h00;
memory3_reg[845 ] <= 8'h00;
memory3_reg[846 ] <= 8'h00;
memory3_reg[847 ] <= 8'h00;
memory3_reg[848 ] <= 8'h00;
memory3_reg[849 ] <= 8'h00;
memory3_reg[850 ] <= 8'h00;
memory3_reg[851 ] <= 8'h00;
memory3_reg[852 ] <= 8'h00;
memory3_reg[853 ] <= 8'h00;
memory3_reg[854 ] <= 8'h00;
memory3_reg[855 ] <= 8'h00;
memory3_reg[856 ] <= 8'h00;
memory3_reg[857 ] <= 8'h00;
memory3_reg[858 ] <= 8'h00;
memory3_reg[859 ] <= 8'h00;
memory3_reg[860 ] <= 8'h00;
memory3_reg[861 ] <= 8'h00;
memory3_reg[862 ] <= 8'h00;
memory3_reg[863 ] <= 8'h00;
memory3_reg[864 ] <= 8'h00;
memory3_reg[865 ] <= 8'h00;
memory3_reg[866 ] <= 8'h00;
memory3_reg[867 ] <= 8'h00;
memory3_reg[868 ] <= 8'h00;
memory3_reg[869 ] <= 8'h00;
memory3_reg[870 ] <= 8'h00;
memory3_reg[871 ] <= 8'h00;
memory3_reg[872 ] <= 8'h00;
memory3_reg[873 ] <= 8'h00;
memory3_reg[874 ] <= 8'h00;
memory3_reg[875 ] <= 8'h00;
memory3_reg[876 ] <= 8'h00;
memory3_reg[877 ] <= 8'h00;
memory3_reg[878 ] <= 8'h00;
memory3_reg[879 ] <= 8'h00;
memory3_reg[880 ] <= 8'h00;
memory3_reg[881 ] <= 8'h00;
memory3_reg[882 ] <= 8'h00;
memory3_reg[883 ] <= 8'h00;
memory3_reg[884 ] <= 8'h00;
memory3_reg[885 ] <= 8'h00;
memory3_reg[886 ] <= 8'h00;
memory3_reg[887 ] <= 8'h00;
memory3_reg[888 ] <= 8'h00;
memory3_reg[889 ] <= 8'h00;
memory3_reg[890 ] <= 8'h00;
memory3_reg[891 ] <= 8'h00;
memory3_reg[892 ] <= 8'h00;
memory3_reg[893 ] <= 8'h00;
memory3_reg[894 ] <= 8'h00;
memory3_reg[895 ] <= 8'h00;
memory3_reg[896 ] <= 8'h00;
memory3_reg[897 ] <= 8'h00;
memory3_reg[898 ] <= 8'h00;
memory3_reg[899 ] <= 8'h00;
memory3_reg[900 ] <= 8'h00;
memory3_reg[901 ] <= 8'h00;
memory3_reg[902 ] <= 8'h00;
memory3_reg[903 ] <= 8'h00;
memory3_reg[904 ] <= 8'h00;
memory3_reg[905 ] <= 8'h00;
memory3_reg[906 ] <= 8'h00;
memory3_reg[907 ] <= 8'h00;
memory3_reg[908 ] <= 8'h00;
memory3_reg[909 ] <= 8'h00;
memory3_reg[910 ] <= 8'h00;
memory3_reg[911 ] <= 8'h00;
memory3_reg[912 ] <= 8'h00;
memory3_reg[913 ] <= 8'h00;
memory3_reg[914 ] <= 8'h00;
memory3_reg[915 ] <= 8'h00;
memory3_reg[916 ] <= 8'h00;
memory3_reg[917 ] <= 8'h00;
memory3_reg[918 ] <= 8'h00;
memory3_reg[919 ] <= 8'h00;
memory3_reg[920 ] <= 8'h00;
memory3_reg[921 ] <= 8'h00;
memory3_reg[922 ] <= 8'h00;
memory3_reg[923 ] <= 8'h00;
memory3_reg[924 ] <= 8'h00;
memory3_reg[925 ] <= 8'h00;
memory3_reg[926 ] <= 8'h00;
memory3_reg[927 ] <= 8'h00;
memory3_reg[928 ] <= 8'h00;
memory3_reg[929 ] <= 8'h00;
memory3_reg[930 ] <= 8'h00;
memory3_reg[931 ] <= 8'h00;
memory3_reg[932 ] <= 8'h00;
memory3_reg[933 ] <= 8'h00;
memory3_reg[934 ] <= 8'h00;
memory3_reg[935 ] <= 8'h00;
memory3_reg[936 ] <= 8'h00;
memory3_reg[937 ] <= 8'h00;
memory3_reg[938 ] <= 8'h00;
memory3_reg[939 ] <= 8'h00;
memory3_reg[940 ] <= 8'h00;
memory3_reg[941 ] <= 8'h00;
memory3_reg[942 ] <= 8'h00;
memory3_reg[943 ] <= 8'h00;
memory3_reg[944 ] <= 8'h00;
memory3_reg[945 ] <= 8'h00;
memory3_reg[946 ] <= 8'h00;
memory3_reg[947 ] <= 8'h00;
memory3_reg[948 ] <= 8'h00;
memory3_reg[949 ] <= 8'h00;
memory3_reg[950 ] <= 8'h00;
memory3_reg[951 ] <= 8'h00;
memory3_reg[952 ] <= 8'h00;
memory3_reg[953 ] <= 8'h00;
memory3_reg[954 ] <= 8'h00;
memory3_reg[955 ] <= 8'h00;
memory3_reg[956 ] <= 8'h00;
memory3_reg[957 ] <= 8'h00;
memory3_reg[958 ] <= 8'h00;
memory3_reg[959 ] <= 8'h00;
memory3_reg[960 ] <= 8'h00;
memory3_reg[961 ] <= 8'h00;
memory3_reg[962 ] <= 8'h00;
memory3_reg[963 ] <= 8'h00;
memory3_reg[964 ] <= 8'h00;
memory3_reg[965 ] <= 8'h00;
memory3_reg[966 ] <= 8'h00;
memory3_reg[967 ] <= 8'h00;
memory3_reg[968 ] <= 8'h00;
memory3_reg[969 ] <= 8'h00;
memory3_reg[970 ] <= 8'h00;
memory3_reg[971 ] <= 8'h00;
memory3_reg[972 ] <= 8'h00;
memory3_reg[973 ] <= 8'h00;
memory3_reg[974 ] <= 8'h00;
memory3_reg[975 ] <= 8'h00;
memory3_reg[976 ] <= 8'h00;
memory3_reg[977 ] <= 8'h00;
memory3_reg[978 ] <= 8'h00;
memory3_reg[979 ] <= 8'h00;
memory3_reg[980 ] <= 8'h00;
memory3_reg[981 ] <= 8'h00;
memory3_reg[982 ] <= 8'h00;
memory3_reg[983 ] <= 8'h00;
memory3_reg[984 ] <= 8'h00;
memory3_reg[985 ] <= 8'h00;
memory3_reg[986 ] <= 8'h00;
memory3_reg[987 ] <= 8'h00;
memory3_reg[988 ] <= 8'h00;
memory3_reg[989 ] <= 8'h00;
memory3_reg[990 ] <= 8'h00;
memory3_reg[991 ] <= 8'h00;
memory3_reg[992 ] <= 8'h00;
memory3_reg[993 ] <= 8'h00;
memory3_reg[994 ] <= 8'h00;
memory3_reg[995 ] <= 8'h00;
memory3_reg[996 ] <= 8'h00;
memory3_reg[997 ] <= 8'h00;
memory3_reg[998 ] <= 8'h00;
memory3_reg[999 ] <= 8'h00;
memory3_reg[1000] <= 8'h00;
memory3_reg[1001] <= 8'h00;
memory3_reg[1002] <= 8'h00;
memory3_reg[1003] <= 8'h00;
memory3_reg[1004] <= 8'h00;
memory3_reg[1005] <= 8'h00;
memory3_reg[1006] <= 8'h00;
memory3_reg[1007] <= 8'h00;
memory3_reg[1008] <= 8'h00;
memory3_reg[1009] <= 8'h00;
memory3_reg[1010] <= 8'h00;
memory3_reg[1011] <= 8'h00;
memory3_reg[1012] <= 8'h00;
memory3_reg[1013] <= 8'h00;
memory3_reg[1014] <= 8'h00;
memory3_reg[1015] <= 8'h00;
memory3_reg[1016] <= 8'h00;
memory3_reg[1017] <= 8'h00;
memory3_reg[1018] <= 8'h00;
memory3_reg[1019] <= 8'h00;
memory3_reg[1020] <= 8'h00;
memory3_reg[1021] <= 8'h00;
memory3_reg[1022] <= 8'h00;
memory3_reg[1023] <= 8'h00;

end

always @(posedge clk_a) begin
    memory0 <= memory0_reg[address_a];
end

always @(posedge clk_a) begin
    memory1 <= memory1_reg[address_a];
end

always @(posedge clk_a) begin
    memory2 <= memory2_reg[address_a];
end

always @(posedge clk_a) begin
    memory3 <= memory3_reg[address_a];
end

assign q_a = {memory0[3:0], memory1[3:0], memory2[3:0], memory3[3:0]};
endmodule