`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.05.2023 09:26:30
// Design Name: 
// Module Name: Sound_program_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CPU_program_rom_2(
    input               clk,
    input       [12:0]  address,
    output reg  [7:0]   data
    );
    
    reg [7:0] ROM_MEM [8191:0];
    integer i;
    initial begin
    ROM_MEM[0   ] <= 8'h08;
ROM_MEM[1   ] <= 8'h38;
ROM_MEM[2   ] <= 8'h00;
ROM_MEM[3   ] <= 8'h20;
ROM_MEM[4   ] <= 8'h00;
ROM_MEM[5   ] <= 8'h01;
ROM_MEM[6   ] <= 8'h00;
ROM_MEM[7   ] <= 8'h09;
ROM_MEM[8   ] <= 8'h38;
ROM_MEM[9   ] <= 8'h00;
ROM_MEM[10  ] <= 8'h50;
ROM_MEM[11  ] <= 8'h00;
ROM_MEM[12  ] <= 8'h01;
ROM_MEM[13  ] <= 8'h03;
ROM_MEM[14  ] <= 8'h0A;
ROM_MEM[15  ] <= 8'h48;
ROM_MEM[16  ] <= 8'h00;
ROM_MEM[17  ] <= 8'hE8;
ROM_MEM[18  ] <= 8'h00;
ROM_MEM[19  ] <= 8'h01;
ROM_MEM[20  ] <= 8'h00;
ROM_MEM[21  ] <= 8'h0B;
ROM_MEM[22  ] <= 8'h48;
ROM_MEM[23  ] <= 8'h00;
ROM_MEM[24  ] <= 8'h18;
ROM_MEM[25  ] <= 8'h00;
ROM_MEM[26  ] <= 8'h01;
ROM_MEM[27  ] <= 8'h00;
ROM_MEM[28  ] <= 8'h0C;
ROM_MEM[29  ] <= 8'h50;
ROM_MEM[30  ] <= 8'h00;
ROM_MEM[31  ] <= 8'h88;
ROM_MEM[32  ] <= 8'h00;
ROM_MEM[33  ] <= 8'h01;
ROM_MEM[34  ] <= 8'h02;
ROM_MEM[35  ] <= 8'h0D;
ROM_MEM[36  ] <= 8'h50;
ROM_MEM[37  ] <= 8'h00;
ROM_MEM[38  ] <= 8'hA0;
ROM_MEM[39  ] <= 8'h00;
ROM_MEM[40  ] <= 8'h01;
ROM_MEM[41  ] <= 8'h03;
ROM_MEM[42  ] <= 8'h0E;
ROM_MEM[43  ] <= 8'h50;
ROM_MEM[44  ] <= 8'h00;
ROM_MEM[45  ] <= 8'hC0;
ROM_MEM[46  ] <= 8'h00;
ROM_MEM[47  ] <= 8'h01;
ROM_MEM[48  ] <= 8'h01;
ROM_MEM[49  ] <= 8'h0F;
ROM_MEM[50  ] <= 8'h50;
ROM_MEM[51  ] <= 8'h00;
ROM_MEM[52  ] <= 8'h40;
ROM_MEM[53  ] <= 8'h00;
ROM_MEM[54  ] <= 8'h01;
ROM_MEM[55  ] <= 8'h01;
ROM_MEM[56  ] <= 8'h10;
ROM_MEM[57  ] <= 8'h50;
ROM_MEM[58  ] <= 8'h00;
ROM_MEM[59  ] <= 8'h60;
ROM_MEM[60  ] <= 8'h00;
ROM_MEM[61  ] <= 8'h01;
ROM_MEM[62  ] <= 8'h03;
ROM_MEM[63  ] <= 8'h11;
ROM_MEM[64  ] <= 8'h50;
ROM_MEM[65  ] <= 8'h00;
ROM_MEM[66  ] <= 8'h78;
ROM_MEM[67  ] <= 8'h00;
ROM_MEM[68  ] <= 8'h01;
ROM_MEM[69  ] <= 8'h02;
ROM_MEM[70  ] <= 8'h12;
ROM_MEM[71  ] <= 8'h5C;
ROM_MEM[72  ] <= 8'h00;
ROM_MEM[73  ] <= 8'hE4;
ROM_MEM[74  ] <= 8'h00;
ROM_MEM[75  ] <= 8'h01;
ROM_MEM[76  ] <= 8'h00;
ROM_MEM[77  ] <= 8'h13;
ROM_MEM[78  ] <= 8'h5C;
ROM_MEM[79  ] <= 8'h00;
ROM_MEM[80  ] <= 8'h1C;
ROM_MEM[81  ] <= 8'h00;
ROM_MEM[82  ] <= 8'h01;
ROM_MEM[83  ] <= 8'h00;
ROM_MEM[84  ] <= 8'h14;
ROM_MEM[85  ] <= 8'h60;
ROM_MEM[86  ] <= 8'h00;
ROM_MEM[87  ] <= 8'hF0;
ROM_MEM[88  ] <= 8'h00;
ROM_MEM[89  ] <= 8'h01;
ROM_MEM[90  ] <= 8'h00;
ROM_MEM[91  ] <= 8'h15;
ROM_MEM[92  ] <= 8'h60;
ROM_MEM[93  ] <= 8'h00;
ROM_MEM[94  ] <= 8'h10;
ROM_MEM[95  ] <= 8'h00;
ROM_MEM[96  ] <= 8'h01;
ROM_MEM[97  ] <= 8'h00;
ROM_MEM[98  ] <= 8'h16;
ROM_MEM[99  ] <= 8'h60;
ROM_MEM[100 ] <= 8'h00;
ROM_MEM[101 ] <= 8'h7C;
ROM_MEM[102 ] <= 8'h00;
ROM_MEM[103 ] <= 8'h01;
ROM_MEM[104 ] <= 8'h03;
ROM_MEM[105 ] <= 8'h17;
ROM_MEM[106 ] <= 8'h70;
ROM_MEM[107 ] <= 8'h00;
ROM_MEM[108 ] <= 8'hC8;
ROM_MEM[109 ] <= 8'h00;
ROM_MEM[110 ] <= 8'h01;
ROM_MEM[111 ] <= 8'h01;
ROM_MEM[112 ] <= 8'h18;
ROM_MEM[113 ] <= 8'h70;
ROM_MEM[114 ] <= 8'h00;
ROM_MEM[115 ] <= 8'hF8;
ROM_MEM[116 ] <= 8'h00;
ROM_MEM[117 ] <= 8'h01;
ROM_MEM[118 ] <= 8'h00;
ROM_MEM[119 ] <= 8'h19;
ROM_MEM[120 ] <= 8'h70;
ROM_MEM[121 ] <= 8'h00;
ROM_MEM[122 ] <= 8'h08;
ROM_MEM[123 ] <= 8'h00;
ROM_MEM[124 ] <= 8'h01;
ROM_MEM[125 ] <= 8'h00;
ROM_MEM[126 ] <= 8'h1A;
ROM_MEM[127 ] <= 8'h70;
ROM_MEM[128 ] <= 8'h00;
ROM_MEM[129 ] <= 8'h38;
ROM_MEM[130 ] <= 8'h00;
ROM_MEM[131 ] <= 8'h01;
ROM_MEM[132 ] <= 8'h01;
ROM_MEM[133 ] <= 8'h1B;
ROM_MEM[134 ] <= 8'h00;
ROM_MEM[135 ] <= 8'h00;
ROM_MEM[136 ] <= 8'hA0;
ROM_MEM[137 ] <= 8'h00;
ROM_MEM[138 ] <= 8'h01;
ROM_MEM[139 ] <= 8'h03;
ROM_MEM[140 ] <= 8'h1C;
ROM_MEM[141 ] <= 8'h00;
ROM_MEM[142 ] <= 8'h00;
ROM_MEM[143 ] <= 8'hC0;
ROM_MEM[144 ] <= 8'h00;
ROM_MEM[145 ] <= 8'h01;
ROM_MEM[146 ] <= 8'h02;
ROM_MEM[147 ] <= 8'h1D;
ROM_MEM[148 ] <= 8'h00;
ROM_MEM[149 ] <= 8'h00;
ROM_MEM[150 ] <= 8'h40;
ROM_MEM[151 ] <= 8'h00;
ROM_MEM[152 ] <= 8'h01;
ROM_MEM[153 ] <= 8'h02;
ROM_MEM[154 ] <= 8'h1E;
ROM_MEM[155 ] <= 8'h00;
ROM_MEM[156 ] <= 8'h00;
ROM_MEM[157 ] <= 8'h60;
ROM_MEM[158 ] <= 8'h00;
ROM_MEM[159 ] <= 8'h01;
ROM_MEM[160 ] <= 8'h03;
ROM_MEM[161 ] <= 8'h1F;
ROM_MEM[162 ] <= 8'h10;
ROM_MEM[163 ] <= 8'h00;
ROM_MEM[164 ] <= 8'hE0;
ROM_MEM[165 ] <= 8'h00;
ROM_MEM[166 ] <= 8'h01;
ROM_MEM[167 ] <= 8'h01;
ROM_MEM[168 ] <= 8'h00;
ROM_MEM[169 ] <= 8'h10;
ROM_MEM[170 ] <= 8'h00;
ROM_MEM[171 ] <= 8'h20;
ROM_MEM[172 ] <= 8'h00;
ROM_MEM[173 ] <= 8'h01;
ROM_MEM[174 ] <= 8'h01;
ROM_MEM[175 ] <= 8'h01;
ROM_MEM[176 ] <= 8'h20;
ROM_MEM[177 ] <= 8'h00;
ROM_MEM[178 ] <= 8'hC0;
ROM_MEM[179 ] <= 8'h00;
ROM_MEM[180 ] <= 8'h03;
ROM_MEM[181 ] <= 8'h01;
ROM_MEM[182 ] <= 8'h02;
ROM_MEM[183 ] <= 8'h20;
ROM_MEM[184 ] <= 8'h00;
ROM_MEM[185 ] <= 8'h40;
ROM_MEM[186 ] <= 8'h00;
ROM_MEM[187 ] <= 8'h03;
ROM_MEM[188 ] <= 8'h01;
ROM_MEM[189 ] <= 8'h03;
ROM_MEM[190 ] <= 8'h28;
ROM_MEM[191 ] <= 8'h00;
ROM_MEM[192 ] <= 8'hE0;
ROM_MEM[193 ] <= 8'h00;
ROM_MEM[194 ] <= 8'h01;
ROM_MEM[195 ] <= 8'h00;
ROM_MEM[196 ] <= 8'h04;
ROM_MEM[197 ] <= 8'h28;
ROM_MEM[198 ] <= 8'h00;
ROM_MEM[199 ] <= 8'h20;
ROM_MEM[200 ] <= 8'h00;
ROM_MEM[201 ] <= 8'h01;
ROM_MEM[202 ] <= 8'h00;
ROM_MEM[203 ] <= 8'h05;
ROM_MEM[204 ] <= 8'h30;
ROM_MEM[205 ] <= 8'h00;
ROM_MEM[206 ] <= 8'h90;
ROM_MEM[207 ] <= 8'h00;
ROM_MEM[208 ] <= 8'h03;
ROM_MEM[209 ] <= 8'h02;
ROM_MEM[210 ] <= 8'h06;
ROM_MEM[211 ] <= 8'h30;
ROM_MEM[212 ] <= 8'h00;
ROM_MEM[213 ] <= 8'hA0;
ROM_MEM[214 ] <= 8'h00;
ROM_MEM[215 ] <= 8'h03;
ROM_MEM[216 ] <= 8'h02;
ROM_MEM[217 ] <= 8'h07;
ROM_MEM[218 ] <= 8'h30;
ROM_MEM[219 ] <= 8'h00;
ROM_MEM[220 ] <= 8'h60;
ROM_MEM[221 ] <= 8'h00;
ROM_MEM[222 ] <= 8'h03;
ROM_MEM[223 ] <= 8'h02;
ROM_MEM[224 ] <= 8'h08;
ROM_MEM[225 ] <= 8'h38;
ROM_MEM[226 ] <= 8'h00;
ROM_MEM[227 ] <= 8'hB0;
ROM_MEM[228 ] <= 8'h00;
ROM_MEM[229 ] <= 8'h01;
ROM_MEM[230 ] <= 8'h01;
ROM_MEM[231 ] <= 8'h09;
ROM_MEM[232 ] <= 8'h38;
ROM_MEM[233 ] <= 8'h00;
ROM_MEM[234 ] <= 8'h50;
ROM_MEM[235 ] <= 8'h00;
ROM_MEM[236 ] <= 8'h01;
ROM_MEM[237 ] <= 8'h01;
ROM_MEM[238 ] <= 8'h0A;
ROM_MEM[239 ] <= 8'h40;
ROM_MEM[240 ] <= 8'h00;
ROM_MEM[241 ] <= 8'hD0;
ROM_MEM[242 ] <= 8'h00;
ROM_MEM[243 ] <= 8'h03;
ROM_MEM[244 ] <= 8'h00;
ROM_MEM[245 ] <= 8'h0B;
ROM_MEM[246 ] <= 8'h40;
ROM_MEM[247 ] <= 8'h00;
ROM_MEM[248 ] <= 8'h00;
ROM_MEM[249 ] <= 8'h00;
ROM_MEM[250 ] <= 8'h03;
ROM_MEM[251 ] <= 8'h00;
ROM_MEM[252 ] <= 8'h0C;
ROM_MEM[253 ] <= 8'h40;
ROM_MEM[254 ] <= 8'h00;
ROM_MEM[255 ] <= 8'h30;
ROM_MEM[256 ] <= 8'h00;
ROM_MEM[257 ] <= 8'h03;
ROM_MEM[258 ] <= 8'h00;
ROM_MEM[259 ] <= 8'h0D;
ROM_MEM[260 ] <= 8'h40;
ROM_MEM[261 ] <= 8'h00;
ROM_MEM[262 ] <= 8'h80;
ROM_MEM[263 ] <= 8'h00;
ROM_MEM[264 ] <= 8'h01;
ROM_MEM[265 ] <= 8'h01;
ROM_MEM[266 ] <= 8'h0E;
ROM_MEM[267 ] <= 8'h50;
ROM_MEM[268 ] <= 8'h00;
ROM_MEM[269 ] <= 8'h88;
ROM_MEM[270 ] <= 8'h00;
ROM_MEM[271 ] <= 8'h01;
ROM_MEM[272 ] <= 8'h02;
ROM_MEM[273 ] <= 8'h0F;
ROM_MEM[274 ] <= 8'h50;
ROM_MEM[275 ] <= 8'h00;
ROM_MEM[276 ] <= 8'h00;
ROM_MEM[277 ] <= 8'h00;
ROM_MEM[278 ] <= 8'h01;
ROM_MEM[279 ] <= 8'h00;
ROM_MEM[280 ] <= 8'h10;
ROM_MEM[281 ] <= 8'h50;
ROM_MEM[282 ] <= 8'h00;
ROM_MEM[283 ] <= 8'h78;
ROM_MEM[284 ] <= 8'h00;
ROM_MEM[285 ] <= 8'h01;
ROM_MEM[286 ] <= 8'h02;
ROM_MEM[287 ] <= 8'h11;
ROM_MEM[288 ] <= 8'h60;
ROM_MEM[289 ] <= 8'h00;
ROM_MEM[290 ] <= 8'hC0;
ROM_MEM[291 ] <= 8'h00;
ROM_MEM[292 ] <= 8'h01;
ROM_MEM[293 ] <= 8'h00;
ROM_MEM[294 ] <= 8'h12;
ROM_MEM[295 ] <= 8'h60;
ROM_MEM[296 ] <= 8'h00;
ROM_MEM[297 ] <= 8'h40;
ROM_MEM[298 ] <= 8'h00;
ROM_MEM[299 ] <= 8'h01;
ROM_MEM[300 ] <= 8'h00;
ROM_MEM[301 ] <= 8'h13;
ROM_MEM[302 ] <= 8'h68;
ROM_MEM[303 ] <= 8'h00;
ROM_MEM[304 ] <= 8'hD0;
ROM_MEM[305 ] <= 8'h00;
ROM_MEM[306 ] <= 8'h01;
ROM_MEM[307 ] <= 8'h00;
ROM_MEM[308 ] <= 8'h14;
ROM_MEM[309 ] <= 8'h68;
ROM_MEM[310 ] <= 8'h00;
ROM_MEM[311 ] <= 8'h30;
ROM_MEM[312 ] <= 8'h00;
ROM_MEM[313 ] <= 8'h01;
ROM_MEM[314 ] <= 8'h00;
ROM_MEM[315 ] <= 8'h15;
ROM_MEM[316 ] <= 8'h70;
ROM_MEM[317 ] <= 8'h00;
ROM_MEM[318 ] <= 8'h90;
ROM_MEM[319 ] <= 8'h00;
ROM_MEM[320 ] <= 8'h01;
ROM_MEM[321 ] <= 8'h01;
ROM_MEM[322 ] <= 8'h16;
ROM_MEM[323 ] <= 8'h70;
ROM_MEM[324 ] <= 8'h00;
ROM_MEM[325 ] <= 8'hA0;
ROM_MEM[326 ] <= 8'h00;
ROM_MEM[327 ] <= 8'h01;
ROM_MEM[328 ] <= 8'h01;
ROM_MEM[329 ] <= 8'h17;
ROM_MEM[330 ] <= 8'h70;
ROM_MEM[331 ] <= 8'h00;
ROM_MEM[332 ] <= 8'hF0;
ROM_MEM[333 ] <= 8'h00;
ROM_MEM[334 ] <= 8'h01;
ROM_MEM[335 ] <= 8'h00;
ROM_MEM[336 ] <= 8'h18;
ROM_MEM[337 ] <= 8'h70;
ROM_MEM[338 ] <= 8'h00;
ROM_MEM[339 ] <= 8'h10;
ROM_MEM[340 ] <= 8'h00;
ROM_MEM[341 ] <= 8'h01;
ROM_MEM[342 ] <= 8'h00;
ROM_MEM[343 ] <= 8'h19;
ROM_MEM[344 ] <= 8'h70;
ROM_MEM[345 ] <= 8'h00;
ROM_MEM[346 ] <= 8'h60;
ROM_MEM[347 ] <= 8'h00;
ROM_MEM[348 ] <= 8'h01;
ROM_MEM[349 ] <= 8'h01;
ROM_MEM[350 ] <= 8'h1A;
ROM_MEM[351 ] <= 8'h70;
ROM_MEM[352 ] <= 8'h00;
ROM_MEM[353 ] <= 8'h70;
ROM_MEM[354 ] <= 8'h00;
ROM_MEM[355 ] <= 8'h01;
ROM_MEM[356 ] <= 8'h01;
ROM_MEM[357 ] <= 8'h1B;
ROM_MEM[358 ] <= 8'h10;
ROM_MEM[359 ] <= 8'h00;
ROM_MEM[360 ] <= 8'hB8;
ROM_MEM[361 ] <= 8'h00;
ROM_MEM[362 ] <= 8'h01;
ROM_MEM[363 ] <= 8'h02;
ROM_MEM[364 ] <= 8'h1C;
ROM_MEM[365 ] <= 8'h10;
ROM_MEM[366 ] <= 8'h00;
ROM_MEM[367 ] <= 8'h58;
ROM_MEM[368 ] <= 8'h00;
ROM_MEM[369 ] <= 8'h01;
ROM_MEM[370 ] <= 8'h02;
ROM_MEM[371 ] <= 8'h1D;
ROM_MEM[372 ] <= 8'h20;
ROM_MEM[373 ] <= 8'h00;
ROM_MEM[374 ] <= 8'h98;
ROM_MEM[375 ] <= 8'h00;
ROM_MEM[376 ] <= 8'h01;
ROM_MEM[377 ] <= 8'h02;
ROM_MEM[378 ] <= 8'h1E;
ROM_MEM[379 ] <= 8'h20;
ROM_MEM[380 ] <= 8'h00;
ROM_MEM[381 ] <= 8'h70;
ROM_MEM[382 ] <= 8'h00;
ROM_MEM[383 ] <= 8'h01;
ROM_MEM[384 ] <= 8'h02;
ROM_MEM[385 ] <= 8'h1F;
ROM_MEM[386 ] <= 8'h9A;
ROM_MEM[387 ] <= 8'h9E;
ROM_MEM[388 ] <= 8'h9B;
ROM_MEM[389 ] <= 8'h62;
ROM_MEM[390 ] <= 8'h9E;
ROM_MEM[391 ] <= 8'hE2;
ROM_MEM[392 ] <= 8'h9F;
ROM_MEM[393 ] <= 8'hA6;
ROM_MEM[394 ] <= 8'h99;
ROM_MEM[395 ] <= 8'hBE;
ROM_MEM[396 ] <= 8'h9A;
ROM_MEM[397 ] <= 8'h82;
ROM_MEM[398 ] <= 8'hA0;
ROM_MEM[399 ] <= 8'hA2;
ROM_MEM[400 ] <= 8'hA1;
ROM_MEM[401 ] <= 8'h66;
ROM_MEM[402 ] <= 8'h9E;
ROM_MEM[403 ] <= 8'h02;
ROM_MEM[404 ] <= 8'h9E;
ROM_MEM[405 ] <= 8'hC6;
ROM_MEM[406 ] <= 8'h98;
ROM_MEM[407 ] <= 8'hDE;
ROM_MEM[408 ] <= 8'h99;
ROM_MEM[409 ] <= 8'hA2;
ROM_MEM[410 ] <= 8'h9D;
ROM_MEM[411 ] <= 8'h22;
ROM_MEM[412 ] <= 8'h9D;
ROM_MEM[413 ] <= 8'hE6;
ROM_MEM[414 ] <= 8'h9C;
ROM_MEM[415 ] <= 8'h42;
ROM_MEM[416 ] <= 8'h9D;
ROM_MEM[417 ] <= 8'h06;
ROM_MEM[418 ] <= 8'h9F;
ROM_MEM[419 ] <= 8'hC2;
ROM_MEM[420 ] <= 8'hA0;
ROM_MEM[421 ] <= 8'h86;
ROM_MEM[422 ] <= 8'h9B;
ROM_MEM[423 ] <= 8'h62;
ROM_MEM[424 ] <= 8'h9C;
ROM_MEM[425 ] <= 8'h26;
ROM_MEM[426 ] <= 8'h9E;
ROM_MEM[427 ] <= 8'hE2;
ROM_MEM[428 ] <= 8'h9F;
ROM_MEM[429 ] <= 8'hC2;
ROM_MEM[430 ] <= 8'h99;
ROM_MEM[431 ] <= 8'hBE;
ROM_MEM[432 ] <= 8'h9A;
ROM_MEM[433 ] <= 8'h9E;
ROM_MEM[434 ] <= 8'hA0;
ROM_MEM[435 ] <= 8'hA2;
ROM_MEM[436 ] <= 8'hA1;
ROM_MEM[437 ] <= 8'h82;
ROM_MEM[438 ] <= 8'h9E;
ROM_MEM[439 ] <= 8'h02;
ROM_MEM[440 ] <= 8'h9E;
ROM_MEM[441 ] <= 8'hE2;
ROM_MEM[442 ] <= 8'h98;
ROM_MEM[443 ] <= 8'hDE;
ROM_MEM[444 ] <= 8'h99;
ROM_MEM[445 ] <= 8'hBE;
ROM_MEM[446 ] <= 8'h9D;
ROM_MEM[447 ] <= 8'h22;
ROM_MEM[448 ] <= 8'h9E;
ROM_MEM[449 ] <= 8'h02;
ROM_MEM[450 ] <= 8'h9C;
ROM_MEM[451 ] <= 8'h42;
ROM_MEM[452 ] <= 8'h9D;
ROM_MEM[453 ] <= 8'h22;
ROM_MEM[454 ] <= 8'h9F;
ROM_MEM[455 ] <= 8'hC2;
ROM_MEM[456 ] <= 8'hA0;
ROM_MEM[457 ] <= 8'hA2;
ROM_MEM[458 ] <= 8'h9B;
ROM_MEM[459 ] <= 8'h62;
ROM_MEM[460 ] <= 8'h9C;
ROM_MEM[461 ] <= 8'h42;
ROM_MEM[462 ] <= 8'hCE;
ROM_MEM[463 ] <= 8'h49;
ROM_MEM[464 ] <= 8'hC2;
ROM_MEM[465 ] <= 8'h86;
ROM_MEM[466 ] <= 8'h00;
ROM_MEM[467 ] <= 8'hA7;
ROM_MEM[468 ] <= 8'hC4;
ROM_MEM[469 ] <= 8'h33;
ROM_MEM[470 ] <= 8'h41;
ROM_MEM[471 ] <= 8'h11;
ROM_MEM[472 ] <= 8'h83;
ROM_MEM[473 ] <= 8'h49;
ROM_MEM[474 ] <= 8'hE2;
ROM_MEM[475 ] <= 8'h25;
ROM_MEM[476 ] <= 8'hF4;
ROM_MEM[477 ] <= 8'hB6;
ROM_MEM[478 ] <= 8'h4B;
ROM_MEM[479 ] <= 8'h13;
ROM_MEM[480 ] <= 8'h81;
ROM_MEM[481 ] <= 8'h13;
ROM_MEM[482 ] <= 8'h25;
ROM_MEM[483 ] <= 8'h0B;
ROM_MEM[484 ] <= 8'hC6;
ROM_MEM[485 ] <= 8'h06;
ROM_MEM[486 ] <= 8'hB6;
ROM_MEM[487 ] <= 8'h47;
ROM_MEM[488 ] <= 8'h03;
ROM_MEM[489 ] <= 8'h3D;
ROM_MEM[490 ] <= 8'h8B;
ROM_MEM[491 ] <= 8'h0D;
ROM_MEM[492 ] <= 8'hB7;
ROM_MEM[493 ] <= 8'h4B;
ROM_MEM[494 ] <= 8'h13;
ROM_MEM[495 ] <= 8'hF6;
ROM_MEM[496 ] <= 8'h4B;
ROM_MEM[497 ] <= 8'h13;
ROM_MEM[498 ] <= 8'h8E;
ROM_MEM[499 ] <= 8'h98;
ROM_MEM[500 ] <= 8'hCB;
ROM_MEM[501 ] <= 8'h3A;
ROM_MEM[502 ] <= 8'h8C;
ROM_MEM[503 ] <= 8'h98;
ROM_MEM[504 ] <= 8'hDE;
ROM_MEM[505 ] <= 8'h25;
ROM_MEM[506 ] <= 8'h03;
ROM_MEM[507 ] <= 8'h8E;
ROM_MEM[508 ] <= 8'h98;
ROM_MEM[509 ] <= 8'hDD;
ROM_MEM[510 ] <= 8'hA6;
ROM_MEM[511 ] <= 8'h84;
ROM_MEM[512 ] <= 8'hB7;
ROM_MEM[513 ] <= 8'h4B;
ROM_MEM[514 ] <= 8'h1A;
ROM_MEM[515 ] <= 8'hFC;
ROM_MEM[516 ] <= 8'h98;
ROM_MEM[517 ] <= 8'h56;
ROM_MEM[518 ] <= 8'hFD;
ROM_MEM[519 ] <= 8'h4B;
ROM_MEM[520 ] <= 8'h2E;
ROM_MEM[521 ] <= 8'hB6;
ROM_MEM[522 ] <= 8'h98;
ROM_MEM[523 ] <= 8'h58;
ROM_MEM[524 ] <= 8'hB7;
ROM_MEM[525 ] <= 8'h4B;
ROM_MEM[526 ] <= 8'h30;
ROM_MEM[527 ] <= 8'h86;
ROM_MEM[528 ] <= 8'h00;
ROM_MEM[529 ] <= 8'h97;
ROM_MEM[530 ] <= 8'hA7;
ROM_MEM[531 ] <= 8'h39;
ROM_MEM[532 ] <= 8'hC6;
ROM_MEM[533 ] <= 8'h07;
ROM_MEM[534 ] <= 8'hD7;
ROM_MEM[535 ] <= 8'hDC;
ROM_MEM[536 ] <= 8'hBD;
ROM_MEM[537 ] <= 8'hCD;
ROM_MEM[538 ] <= 8'h38;
ROM_MEM[539 ] <= 8'hCC;
ROM_MEM[540 ] <= 8'h00;
ROM_MEM[541 ] <= 8'h00;
ROM_MEM[542 ] <= 8'hFD;
ROM_MEM[543 ] <= 8'h50;
ROM_MEM[544 ] <= 8'h40;
ROM_MEM[545 ] <= 8'hFD;
ROM_MEM[546 ] <= 8'h50;
ROM_MEM[547 ] <= 8'h42;
ROM_MEM[548 ] <= 8'hFD;
ROM_MEM[549 ] <= 8'h50;
ROM_MEM[550 ] <= 8'h44;
ROM_MEM[551 ] <= 8'hBD;
ROM_MEM[552 ] <= 8'hA4;
ROM_MEM[553 ] <= 8'h0A;
ROM_MEM[554 ] <= 8'hFC;
ROM_MEM[555 ] <= 8'h50;
ROM_MEM[556 ] <= 8'h98;
ROM_MEM[557 ] <= 8'hFD;
ROM_MEM[558 ] <= 8'h50;
ROM_MEM[559 ] <= 8'h40;
ROM_MEM[560 ] <= 8'hFC;
ROM_MEM[561 ] <= 8'h50;
ROM_MEM[562 ] <= 8'h9A;
ROM_MEM[563 ] <= 8'hFD;
ROM_MEM[564 ] <= 8'h50;
ROM_MEM[565 ] <= 8'h42;
ROM_MEM[566 ] <= 8'hFC;
ROM_MEM[567 ] <= 8'h50;
ROM_MEM[568 ] <= 8'h9C;
ROM_MEM[569 ] <= 8'hFD;
ROM_MEM[570 ] <= 8'h50;
ROM_MEM[571 ] <= 8'h44;
ROM_MEM[572 ] <= 8'hF6;
ROM_MEM[573 ] <= 8'h4B;
ROM_MEM[574 ] <= 8'h13;
ROM_MEM[575 ] <= 8'h58;
ROM_MEM[576 ] <= 8'h58;
ROM_MEM[577 ] <= 8'h8E;
ROM_MEM[578 ] <= 8'hA1;
ROM_MEM[579 ] <= 8'h82;
ROM_MEM[580 ] <= 8'h3A;
ROM_MEM[581 ] <= 8'h8C;
ROM_MEM[582 ] <= 8'hA1;
ROM_MEM[583 ] <= 8'hCE;
ROM_MEM[584 ] <= 8'h25;
ROM_MEM[585 ] <= 8'h03;
ROM_MEM[586 ] <= 8'h8E;
ROM_MEM[587 ] <= 8'hA1;
ROM_MEM[588 ] <= 8'hCA;
ROM_MEM[589 ] <= 8'hAE;
ROM_MEM[590 ] <= 8'h84;
ROM_MEM[591 ] <= 8'h9F;
ROM_MEM[592 ] <= 8'h64;
ROM_MEM[593 ] <= 8'h96;
ROM_MEM[594 ] <= 8'hA7;
ROM_MEM[595 ] <= 8'hA1;
ROM_MEM[596 ] <= 8'h05;
ROM_MEM[597 ] <= 8'h10;
ROM_MEM[598 ] <= 8'h2D;
ROM_MEM[599 ] <= 8'h00;
ROM_MEM[600 ] <= 8'h81;
ROM_MEM[601 ] <= 8'hEC;
ROM_MEM[602 ] <= 8'h84;
ROM_MEM[603 ] <= 8'hFD;
ROM_MEM[604 ] <= 8'h5E;
ROM_MEM[605 ] <= 8'h00;
ROM_MEM[606 ] <= 8'hEC;
ROM_MEM[607 ] <= 8'h02;
ROM_MEM[608 ] <= 8'hFD;
ROM_MEM[609 ] <= 8'h5E;
ROM_MEM[610 ] <= 8'h02;
ROM_MEM[611 ] <= 8'hCC;
ROM_MEM[612 ] <= 8'h1E;
ROM_MEM[613 ] <= 8'h00;
ROM_MEM[614 ] <= 8'hFD;
ROM_MEM[615 ] <= 8'h5E;
ROM_MEM[616 ] <= 8'h04;
ROM_MEM[617 ] <= 8'hCC;
ROM_MEM[618 ] <= 8'h01;
ROM_MEM[619 ] <= 8'hC0;
ROM_MEM[620 ] <= 8'hFD;
ROM_MEM[621 ] <= 8'h47;
ROM_MEM[622 ] <= 8'h01;
ROM_MEM[623 ] <= 8'h86;
ROM_MEM[624 ] <= 8'h67;
ROM_MEM[625 ] <= 8'hBD;
ROM_MEM[626 ] <= 8'hCD;
ROM_MEM[627 ] <= 8'hBA;
ROM_MEM[628 ] <= 8'hFC;
ROM_MEM[629 ] <= 8'h50;
ROM_MEM[630 ] <= 8'h00;
ROM_MEM[631 ] <= 8'h2A;
ROM_MEM[632 ] <= 8'h05;
ROM_MEM[633 ] <= 8'h84;
ROM_MEM[634 ] <= 8'h3F;
ROM_MEM[635 ] <= 8'hFD;
ROM_MEM[636 ] <= 8'h50;
ROM_MEM[637 ] <= 8'h00;
ROM_MEM[638 ] <= 8'hFD;
ROM_MEM[639 ] <= 8'h50;
ROM_MEM[640 ] <= 8'h7C;
ROM_MEM[641 ] <= 8'h10;
ROM_MEM[642 ] <= 8'h83;
ROM_MEM[643 ] <= 8'h01;
ROM_MEM[644 ] <= 8'h00;
ROM_MEM[645 ] <= 8'h2D;
ROM_MEM[646 ] <= 8'h29;
ROM_MEM[647 ] <= 8'h10;
ROM_MEM[648 ] <= 8'h83;
ROM_MEM[649 ] <= 8'h3C;
ROM_MEM[650 ] <= 8'h00;
ROM_MEM[651 ] <= 8'h24;
ROM_MEM[652 ] <= 8'h23;
ROM_MEM[653 ] <= 8'hFC;
ROM_MEM[654 ] <= 8'h50;
ROM_MEM[655 ] <= 8'h02;
ROM_MEM[656 ] <= 8'h2A;
ROM_MEM[657 ] <= 8'h04;
ROM_MEM[658 ] <= 8'h43;
ROM_MEM[659 ] <= 8'h50;
ROM_MEM[660 ] <= 8'h82;
ROM_MEM[661 ] <= 8'hFF;
ROM_MEM[662 ] <= 8'hB3;
ROM_MEM[663 ] <= 8'h50;
ROM_MEM[664 ] <= 8'h00;
ROM_MEM[665 ] <= 8'h24;
ROM_MEM[666 ] <= 8'h15;
ROM_MEM[667 ] <= 8'hCE;
ROM_MEM[668 ] <= 8'h49;
ROM_MEM[669 ] <= 8'hC2;
ROM_MEM[670 ] <= 8'hE6;
ROM_MEM[671 ] <= 8'h06;
ROM_MEM[672 ] <= 8'h33;
ROM_MEM[673 ] <= 8'hC5;
ROM_MEM[674 ] <= 8'hA6;
ROM_MEM[675 ] <= 8'hC4;
ROM_MEM[676 ] <= 8'h85;
ROM_MEM[677 ] <= 8'h02;
ROM_MEM[678 ] <= 8'h27;
ROM_MEM[679 ] <= 8'h06;
ROM_MEM[680 ] <= 8'hBD;
ROM_MEM[681 ] <= 8'hA2;
ROM_MEM[682 ] <= 8'hF8;
ROM_MEM[683 ] <= 8'hBD;
ROM_MEM[684 ] <= 8'hA5;
ROM_MEM[685 ] <= 8'h91;
ROM_MEM[686 ] <= 8'h20;
ROM_MEM[687 ] <= 8'h2A;
ROM_MEM[688 ] <= 8'h9E;
ROM_MEM[689 ] <= 8'h64;
ROM_MEM[690 ] <= 8'hCE;
ROM_MEM[691 ] <= 8'h49;
ROM_MEM[692 ] <= 8'hC2;
ROM_MEM[693 ] <= 8'hE6;
ROM_MEM[694 ] <= 8'h06;
ROM_MEM[695 ] <= 8'h33;
ROM_MEM[696 ] <= 8'hC5;
ROM_MEM[697 ] <= 8'hB6;
ROM_MEM[698 ] <= 8'h4B;
ROM_MEM[699 ] <= 8'h3D;
ROM_MEM[700 ] <= 8'h27;
ROM_MEM[701 ] <= 8'h04;
ROM_MEM[702 ] <= 8'h6F;
ROM_MEM[703 ] <= 8'hC4;
ROM_MEM[704 ] <= 8'h20;
ROM_MEM[705 ] <= 8'h18;
ROM_MEM[706 ] <= 8'h86;
ROM_MEM[707 ] <= 8'h0B;
ROM_MEM[708 ] <= 8'hE6;
ROM_MEM[709 ] <= 8'hC4;
ROM_MEM[710 ] <= 8'hC5;
ROM_MEM[711 ] <= 8'h04;
ROM_MEM[712 ] <= 8'h27;
ROM_MEM[713 ] <= 8'h0C;
ROM_MEM[714 ] <= 8'h8A;
ROM_MEM[715 ] <= 8'h04;
ROM_MEM[716 ] <= 8'hE6;
ROM_MEM[717 ] <= 8'h04;
ROM_MEM[718 ] <= 8'hC1;
ROM_MEM[719 ] <= 8'h03;
ROM_MEM[720 ] <= 8'h26;
ROM_MEM[721 ] <= 8'h02;
ROM_MEM[722 ] <= 8'h84;
ROM_MEM[723 ] <= 8'hFD;
ROM_MEM[724 ] <= 8'h20;
ROM_MEM[725 ] <= 8'h02;
ROM_MEM[726 ] <= 8'h8A;
ROM_MEM[727 ] <= 8'h10;
ROM_MEM[728 ] <= 8'hA7;
ROM_MEM[729 ] <= 8'hC4;
ROM_MEM[730 ] <= 8'hF6;
ROM_MEM[731 ] <= 8'h4B;
ROM_MEM[732 ] <= 8'h13;
ROM_MEM[733 ] <= 8'h58;
ROM_MEM[734 ] <= 8'h58;
ROM_MEM[735 ] <= 8'h8E;
ROM_MEM[736 ] <= 8'hA1;
ROM_MEM[737 ] <= 8'h82;
ROM_MEM[738 ] <= 8'h3A;
ROM_MEM[739 ] <= 8'h8C;
ROM_MEM[740 ] <= 8'hA1;
ROM_MEM[741 ] <= 8'hCE;
ROM_MEM[742 ] <= 8'h25;
ROM_MEM[743 ] <= 8'h03;
ROM_MEM[744 ] <= 8'h8E;
ROM_MEM[745 ] <= 8'hA1;
ROM_MEM[746 ] <= 8'hCA;
ROM_MEM[747 ] <= 8'h1F;
ROM_MEM[748 ] <= 8'h13;
ROM_MEM[749 ] <= 8'h9E;
ROM_MEM[750 ] <= 8'h64;
ROM_MEM[751 ] <= 8'h30;
ROM_MEM[752 ] <= 8'h07;
ROM_MEM[753 ] <= 8'hAC;
ROM_MEM[754 ] <= 8'h42;
ROM_MEM[755 ] <= 8'h10;
ROM_MEM[756 ] <= 8'h25;
ROM_MEM[757 ] <= 8'hFF;
ROM_MEM[758 ] <= 8'h58;
ROM_MEM[759 ] <= 8'h39;
ROM_MEM[760 ] <= 8'h9E;
ROM_MEM[761 ] <= 8'h64;
ROM_MEM[762 ] <= 8'hE6;
ROM_MEM[763 ] <= 8'h04;
ROM_MEM[764 ] <= 8'hC1;
ROM_MEM[765 ] <= 8'h03;
ROM_MEM[766 ] <= 8'h26;
ROM_MEM[767 ] <= 8'h04;
ROM_MEM[768 ] <= 8'hC6;
ROM_MEM[769 ] <= 8'h09;
ROM_MEM[770 ] <= 8'h20;
ROM_MEM[771 ] <= 8'h02;
ROM_MEM[772 ] <= 8'hC6;
ROM_MEM[773 ] <= 8'h08;
ROM_MEM[774 ] <= 8'hD7;
ROM_MEM[775 ] <= 8'hDC;
ROM_MEM[776 ] <= 8'hCC;
ROM_MEM[777 ] <= 8'h66;
ROM_MEM[778 ] <= 8'h80;
ROM_MEM[779 ] <= 8'hFD;
ROM_MEM[780 ] <= 8'h5E;
ROM_MEM[781 ] <= 8'h02;
ROM_MEM[782 ] <= 8'hCE;
ROM_MEM[783 ] <= 8'h49;
ROM_MEM[784 ] <= 8'hC2;
ROM_MEM[785 ] <= 8'hE6;
ROM_MEM[786 ] <= 8'h06;
ROM_MEM[787 ] <= 8'h33;
ROM_MEM[788 ] <= 8'hC5;
ROM_MEM[789 ] <= 8'hA6;
ROM_MEM[790 ] <= 8'hC4;
ROM_MEM[791 ] <= 8'hE6;
ROM_MEM[792 ] <= 8'h04;
ROM_MEM[793 ] <= 8'hC1;
ROM_MEM[794 ] <= 8'h03;
ROM_MEM[795 ] <= 8'h27;
ROM_MEM[796 ] <= 8'h16;
ROM_MEM[797 ] <= 8'h85;
ROM_MEM[798 ] <= 8'h04;
ROM_MEM[799 ] <= 8'h26;
ROM_MEM[800 ] <= 8'h04;
ROM_MEM[801 ] <= 8'h85;
ROM_MEM[802 ] <= 8'h10;
ROM_MEM[803 ] <= 8'h26;
ROM_MEM[804 ] <= 8'h09;
ROM_MEM[805 ] <= 8'hC6;
ROM_MEM[806 ] <= 8'h0A;
ROM_MEM[807 ] <= 8'hD7;
ROM_MEM[808 ] <= 8'hDC;
ROM_MEM[809 ] <= 8'hCC;
ROM_MEM[810 ] <= 8'h60;
ROM_MEM[811 ] <= 8'h80;
ROM_MEM[812 ] <= 8'h20;
ROM_MEM[813 ] <= 8'h03;
ROM_MEM[814 ] <= 8'hCC;
ROM_MEM[815 ] <= 8'h67;
ROM_MEM[816 ] <= 8'h80;
ROM_MEM[817 ] <= 8'h20;
ROM_MEM[818 ] <= 8'h0C;
ROM_MEM[819 ] <= 8'h85;
ROM_MEM[820 ] <= 8'h04;
ROM_MEM[821 ] <= 8'h26;
ROM_MEM[822 ] <= 8'h05;
ROM_MEM[823 ] <= 8'hCC;
ROM_MEM[824 ] <= 8'h64;
ROM_MEM[825 ] <= 8'h60;
ROM_MEM[826 ] <= 8'h20;
ROM_MEM[827 ] <= 8'h03;
ROM_MEM[828 ] <= 8'hCC;
ROM_MEM[829 ] <= 8'h60;
ROM_MEM[830 ] <= 8'h80;
ROM_MEM[831 ] <= 8'hFD;
ROM_MEM[832 ] <= 8'h5E;
ROM_MEM[833 ] <= 8'h00;
ROM_MEM[834 ] <= 8'h86;
ROM_MEM[835 ] <= 8'h72;
ROM_MEM[836 ] <= 8'hB7;
ROM_MEM[837 ] <= 8'h5E;
ROM_MEM[838 ] <= 8'h04;
ROM_MEM[839 ] <= 8'hB6;
ROM_MEM[840 ] <= 8'h50;
ROM_MEM[841 ] <= 8'h00;
ROM_MEM[842 ] <= 8'h48;
ROM_MEM[843 ] <= 8'h48;
ROM_MEM[844 ] <= 8'hB7;
ROM_MEM[845 ] <= 8'h5E;
ROM_MEM[846 ] <= 8'h05;
ROM_MEM[847 ] <= 8'hC6;
ROM_MEM[848 ] <= 8'h40;
ROM_MEM[849 ] <= 8'h43;
ROM_MEM[850 ] <= 8'h3D;
ROM_MEM[851 ] <= 8'h8B;
ROM_MEM[852 ] <= 8'h40;
ROM_MEM[853 ] <= 8'hB7;
ROM_MEM[854 ] <= 8'h5E;
ROM_MEM[855 ] <= 8'h03;
ROM_MEM[856 ] <= 8'hFC;
ROM_MEM[857 ] <= 8'h50;
ROM_MEM[858 ] <= 8'h86;
ROM_MEM[859 ] <= 8'h58;
ROM_MEM[860 ] <= 8'h49;
ROM_MEM[861 ] <= 8'hC3;
ROM_MEM[862 ] <= 8'h04;
ROM_MEM[863 ] <= 8'h00;
ROM_MEM[864 ] <= 8'hB3;
ROM_MEM[865 ] <= 8'h50;
ROM_MEM[866 ] <= 8'h00;
ROM_MEM[867 ] <= 8'h10;
ROM_MEM[868 ] <= 8'h2D;
ROM_MEM[869 ] <= 8'h00;
ROM_MEM[870 ] <= 8'h8D;
ROM_MEM[871 ] <= 8'hA6;
ROM_MEM[872 ] <= 8'h04;
ROM_MEM[873 ] <= 8'h81;
ROM_MEM[874 ] <= 8'h03;
ROM_MEM[875 ] <= 8'h27;
ROM_MEM[876 ] <= 8'h3A;
ROM_MEM[877 ] <= 8'h96;
ROM_MEM[878 ] <= 8'h60;
ROM_MEM[879 ] <= 8'h2D;
ROM_MEM[880 ] <= 8'h03;
ROM_MEM[881 ] <= 8'hBD;
ROM_MEM[882 ] <= 8'hBD;
ROM_MEM[883 ] <= 8'hD0;
ROM_MEM[884 ] <= 8'hFC;
ROM_MEM[885 ] <= 8'h50;
ROM_MEM[886 ] <= 8'h00;
ROM_MEM[887 ] <= 8'h83;
ROM_MEM[888 ] <= 8'h02;
ROM_MEM[889 ] <= 8'h00;
ROM_MEM[890 ] <= 8'hB3;
ROM_MEM[891 ] <= 8'h50;
ROM_MEM[892 ] <= 8'h86;
ROM_MEM[893 ] <= 8'h2E;
ROM_MEM[894 ] <= 8'h26;
ROM_MEM[895 ] <= 8'hCC;
ROM_MEM[896 ] <= 8'hA0;
ROM_MEM[897 ] <= 8'h18;
ROM_MEM[898 ] <= 8'hFD;
ROM_MEM[899 ] <= 8'h5E;
ROM_MEM[900 ] <= 8'h02;
ROM_MEM[901 ] <= 8'hCC;
ROM_MEM[902 ] <= 8'h60;
ROM_MEM[903 ] <= 8'h80;
ROM_MEM[904 ] <= 8'hFD;
ROM_MEM[905 ] <= 8'h5E;
ROM_MEM[906 ] <= 8'h00;
ROM_MEM[907 ] <= 8'h96;
ROM_MEM[908 ] <= 8'h60;
ROM_MEM[909 ] <= 8'h2D;
ROM_MEM[910 ] <= 8'h06;
ROM_MEM[911 ] <= 8'hBD;
ROM_MEM[912 ] <= 8'h98;
ROM_MEM[913 ] <= 8'h74;
ROM_MEM[914 ] <= 8'hBD;
ROM_MEM[915 ] <= 8'hBD;
ROM_MEM[916 ] <= 8'hB2;
ROM_MEM[917 ] <= 8'h96;
ROM_MEM[918 ] <= 8'h63;
ROM_MEM[919 ] <= 8'h26;
ROM_MEM[920 ] <= 8'h04;
ROM_MEM[921 ] <= 8'hB6;
ROM_MEM[922 ] <= 8'h50;
ROM_MEM[923 ] <= 8'h02;
ROM_MEM[924 ] <= 8'h40;
ROM_MEM[925 ] <= 8'hC6;
ROM_MEM[926 ] <= 8'h20;
ROM_MEM[927 ] <= 8'h4D;
ROM_MEM[928 ] <= 8'h2A;
ROM_MEM[929 ] <= 8'h01;
ROM_MEM[930 ] <= 8'h50;
ROM_MEM[931 ] <= 8'hD7;
ROM_MEM[932 ] <= 8'h63;
ROM_MEM[933 ] <= 8'h20;
ROM_MEM[934 ] <= 8'h4D;
ROM_MEM[935 ] <= 8'hFC;
ROM_MEM[936 ] <= 8'h50;
ROM_MEM[937 ] <= 8'h44;
ROM_MEM[938 ] <= 8'h83;
ROM_MEM[939 ] <= 8'h07;
ROM_MEM[940 ] <= 8'hA0;
ROM_MEM[941 ] <= 8'h2E;
ROM_MEM[942 ] <= 8'h45;
ROM_MEM[943 ] <= 8'hBD;
ROM_MEM[944 ] <= 8'hBD;
ROM_MEM[945 ] <= 8'hD0;
ROM_MEM[946 ] <= 8'h9E;
ROM_MEM[947 ] <= 8'h64;
ROM_MEM[948 ] <= 8'hCE;
ROM_MEM[949 ] <= 8'h49;
ROM_MEM[950 ] <= 8'hC2;
ROM_MEM[951 ] <= 8'hE6;
ROM_MEM[952 ] <= 8'h06;
ROM_MEM[953 ] <= 8'h33;
ROM_MEM[954 ] <= 8'hC5;
ROM_MEM[955 ] <= 8'hA6;
ROM_MEM[956 ] <= 8'hC4;
ROM_MEM[957 ] <= 8'h85;
ROM_MEM[958 ] <= 8'h04;
ROM_MEM[959 ] <= 8'h26;
ROM_MEM[960 ] <= 8'h33;
ROM_MEM[961 ] <= 8'hFC;
ROM_MEM[962 ] <= 8'h50;
ROM_MEM[963 ] <= 8'h44;
ROM_MEM[964 ] <= 8'h83;
ROM_MEM[965 ] <= 8'h05;
ROM_MEM[966 ] <= 8'hA0;
ROM_MEM[967 ] <= 8'h2C;
ROM_MEM[968 ] <= 8'h2B;
ROM_MEM[969 ] <= 8'hFC;
ROM_MEM[970 ] <= 8'h50;
ROM_MEM[971 ] <= 8'h00;
ROM_MEM[972 ] <= 8'h83;
ROM_MEM[973 ] <= 8'h04;
ROM_MEM[974 ] <= 8'h00;
ROM_MEM[975 ] <= 8'hB3;
ROM_MEM[976 ] <= 8'h50;
ROM_MEM[977 ] <= 8'h86;
ROM_MEM[978 ] <= 8'h2E;
ROM_MEM[979 ] <= 8'h20;
ROM_MEM[980 ] <= 8'hCC;
ROM_MEM[981 ] <= 8'hA0;
ROM_MEM[982 ] <= 8'h18;
ROM_MEM[983 ] <= 8'hFD;
ROM_MEM[984 ] <= 8'h5E;
ROM_MEM[985 ] <= 8'h00;
ROM_MEM[986 ] <= 8'h96;
ROM_MEM[987 ] <= 8'h60;
ROM_MEM[988 ] <= 8'h2D;
ROM_MEM[989 ] <= 8'h06;
ROM_MEM[990 ] <= 8'hBD;
ROM_MEM[991 ] <= 8'h98;
ROM_MEM[992 ] <= 8'h74;
ROM_MEM[993 ] <= 8'hBD;
ROM_MEM[994 ] <= 8'hBD;
ROM_MEM[995 ] <= 8'hB2;
ROM_MEM[996 ] <= 8'h96;
ROM_MEM[997 ] <= 8'h63;
ROM_MEM[998 ] <= 8'h26;
ROM_MEM[999 ] <= 8'h0C;
ROM_MEM[1000] <= 8'h86;
ROM_MEM[1001] <= 8'h13;
ROM_MEM[1002] <= 8'hF6;
ROM_MEM[1003] <= 8'h50;
ROM_MEM[1004] <= 8'h02;
ROM_MEM[1005] <= 8'h2B;
ROM_MEM[1006] <= 8'h01;
ROM_MEM[1007] <= 8'h40;
ROM_MEM[1008] <= 8'h9B;
ROM_MEM[1009] <= 8'h63;
ROM_MEM[1010] <= 8'h97;
ROM_MEM[1011] <= 8'h63;
ROM_MEM[1012] <= 8'hB6;
ROM_MEM[1013] <= 8'h50;
ROM_MEM[1014] <= 8'h00;
ROM_MEM[1015] <= 8'h80;
ROM_MEM[1016] <= 8'h08;
ROM_MEM[1017] <= 8'h2E;
ROM_MEM[1018] <= 8'h05;
ROM_MEM[1019] <= 8'hBD;
ROM_MEM[1020] <= 8'hCD;
ROM_MEM[1021] <= 8'h68;
ROM_MEM[1022] <= 8'h20;
ROM_MEM[1023] <= 8'h03;
ROM_MEM[1024] <= 8'hBD;
ROM_MEM[1025] <= 8'hCD;
ROM_MEM[1026] <= 8'h50;
ROM_MEM[1027] <= 8'hBD;
ROM_MEM[1028] <= 8'hCD;
ROM_MEM[1029] <= 8'h74;
ROM_MEM[1030] <= 8'hBD;
ROM_MEM[1031] <= 8'hA4;
ROM_MEM[1032] <= 8'h59;
ROM_MEM[1033] <= 8'h39;
ROM_MEM[1034] <= 8'hBD;
ROM_MEM[1035] <= 8'hCD;
ROM_MEM[1036] <= 8'hE7;
ROM_MEM[1037] <= 8'hCC;
ROM_MEM[1038] <= 8'h00;
ROM_MEM[1039] <= 8'h00;
ROM_MEM[1040] <= 8'hFD;
ROM_MEM[1041] <= 8'h50;
ROM_MEM[1042] <= 8'h78;
ROM_MEM[1043] <= 8'hDC;
ROM_MEM[1044] <= 8'hB3;
ROM_MEM[1045] <= 8'hFD;
ROM_MEM[1046] <= 8'h50;
ROM_MEM[1047] <= 8'h7A;
ROM_MEM[1048] <= 8'hDC;
ROM_MEM[1049] <= 8'hB5;
ROM_MEM[1050] <= 8'hFD;
ROM_MEM[1051] <= 8'h50;
ROM_MEM[1052] <= 8'h7C;
ROM_MEM[1053] <= 8'hCC;
ROM_MEM[1054] <= 8'h00;
ROM_MEM[1055] <= 8'h0F;
ROM_MEM[1056] <= 8'hFD;
ROM_MEM[1057] <= 8'h47;
ROM_MEM[1058] <= 8'h01;
ROM_MEM[1059] <= 8'h86;
ROM_MEM[1060] <= 8'h2A;
ROM_MEM[1061] <= 8'hBD;
ROM_MEM[1062] <= 8'hCD;
ROM_MEM[1063] <= 8'hBA;
ROM_MEM[1064] <= 8'hFC;
ROM_MEM[1065] <= 8'h50;
ROM_MEM[1066] <= 8'h02;
ROM_MEM[1067] <= 8'hFD;
ROM_MEM[1068] <= 8'h50;
ROM_MEM[1069] <= 8'h78;
ROM_MEM[1070] <= 8'hFC;
ROM_MEM[1071] <= 8'h50;
ROM_MEM[1072] <= 8'h04;
ROM_MEM[1073] <= 8'hFD;
ROM_MEM[1074] <= 8'h50;
ROM_MEM[1075] <= 8'h7A;
ROM_MEM[1076] <= 8'h2A;
ROM_MEM[1077] <= 8'h1F;
ROM_MEM[1078] <= 8'h96;
ROM_MEM[1079] <= 8'hBC;
ROM_MEM[1080] <= 8'h27;
ROM_MEM[1081] <= 8'h1B;
ROM_MEM[1082] <= 8'h86;
ROM_MEM[1083] <= 8'hFF;
ROM_MEM[1084] <= 8'h97;
ROM_MEM[1085] <= 8'hBD;
ROM_MEM[1086] <= 8'h86;
ROM_MEM[1087] <= 8'h03;
ROM_MEM[1088] <= 8'hB7;
ROM_MEM[1089] <= 8'h4B;
ROM_MEM[1090] <= 8'h23;
ROM_MEM[1091] <= 8'hCC;
ROM_MEM[1092] <= 8'h62;
ROM_MEM[1093] <= 8'h80;
ROM_MEM[1094] <= 8'hFD;
ROM_MEM[1095] <= 8'h4B;
ROM_MEM[1096] <= 8'h20;
ROM_MEM[1097] <= 8'hFC;
ROM_MEM[1098] <= 8'h50;
ROM_MEM[1099] <= 8'h04;
ROM_MEM[1100] <= 8'h44;
ROM_MEM[1101] <= 8'h56;
ROM_MEM[1102] <= 8'h44;
ROM_MEM[1103] <= 8'h56;
ROM_MEM[1104] <= 8'hCB;
ROM_MEM[1105] <= 8'hC0;
ROM_MEM[1106] <= 8'hF7;
ROM_MEM[1107] <= 8'h4B;
ROM_MEM[1108] <= 8'h22;
ROM_MEM[1109] <= 8'hBD;
ROM_MEM[1110] <= 8'hCD;
ROM_MEM[1111] <= 8'hE7;
ROM_MEM[1112] <= 8'h39;
ROM_MEM[1113] <= 8'h9E;
ROM_MEM[1114] <= 8'h64;
ROM_MEM[1115] <= 8'hFC;
ROM_MEM[1116] <= 8'h50;
ROM_MEM[1117] <= 8'h7C;
ROM_MEM[1118] <= 8'h58;
ROM_MEM[1119] <= 8'h49;
ROM_MEM[1120] <= 8'hFD;
ROM_MEM[1121] <= 8'h47;
ROM_MEM[1122] <= 8'h04;
ROM_MEM[1123] <= 8'hEC;
ROM_MEM[1124] <= 8'h02;
ROM_MEM[1125] <= 8'hB3;
ROM_MEM[1126] <= 8'h50;
ROM_MEM[1127] <= 8'h42;
ROM_MEM[1128] <= 8'hFD;
ROM_MEM[1129] <= 8'h50;
ROM_MEM[1130] <= 8'h02;
ROM_MEM[1131] <= 8'hCC;
ROM_MEM[1132] <= 8'h00;
ROM_MEM[1133] <= 8'h00;
ROM_MEM[1134] <= 8'hB3;
ROM_MEM[1135] <= 8'h50;
ROM_MEM[1136] <= 8'h44;
ROM_MEM[1137] <= 8'hFD;
ROM_MEM[1138] <= 8'h50;
ROM_MEM[1139] <= 8'h04;
ROM_MEM[1140] <= 8'hFC;
ROM_MEM[1141] <= 8'h47;
ROM_MEM[1142] <= 8'h00;
ROM_MEM[1143] <= 8'hFD;
ROM_MEM[1144] <= 8'h50;
ROM_MEM[1145] <= 8'h00;
ROM_MEM[1146] <= 8'h86;
ROM_MEM[1147] <= 8'h86;
ROM_MEM[1148] <= 8'hBD;
ROM_MEM[1149] <= 8'hCD;
ROM_MEM[1150] <= 8'hBA;
ROM_MEM[1151] <= 8'hFC;
ROM_MEM[1152] <= 8'h50;
ROM_MEM[1153] <= 8'h02;
ROM_MEM[1154] <= 8'hFD;
ROM_MEM[1155] <= 8'h50;
ROM_MEM[1156] <= 8'h1A;
ROM_MEM[1157] <= 8'hFC;
ROM_MEM[1158] <= 8'h50;
ROM_MEM[1159] <= 8'h04;
ROM_MEM[1160] <= 8'hFD;
ROM_MEM[1161] <= 8'h50;
ROM_MEM[1162] <= 8'h1C;
ROM_MEM[1163] <= 8'hA6;
ROM_MEM[1164] <= 8'h04;
ROM_MEM[1165] <= 8'h81;
ROM_MEM[1166] <= 8'h03;
ROM_MEM[1167] <= 8'h27;
ROM_MEM[1168] <= 8'h0E;
ROM_MEM[1169] <= 8'hCC;
ROM_MEM[1170] <= 8'h03;
ROM_MEM[1171] <= 8'hC0;
ROM_MEM[1172] <= 8'hFD;
ROM_MEM[1173] <= 8'h50;
ROM_MEM[1174] <= 8'h02;
ROM_MEM[1175] <= 8'hCC;
ROM_MEM[1176] <= 8'h52;
ROM_MEM[1177] <= 8'h80;
ROM_MEM[1178] <= 8'hFD;
ROM_MEM[1179] <= 8'h50;
ROM_MEM[1180] <= 8'h04;
ROM_MEM[1181] <= 8'h20;
ROM_MEM[1182] <= 8'h1B;
ROM_MEM[1183] <= 8'hCE;
ROM_MEM[1184] <= 8'h49;
ROM_MEM[1185] <= 8'hC2;
ROM_MEM[1186] <= 8'hE6;
ROM_MEM[1187] <= 8'h06;
ROM_MEM[1188] <= 8'h33;
ROM_MEM[1189] <= 8'hC5;
ROM_MEM[1190] <= 8'hA6;
ROM_MEM[1191] <= 8'hC4;
ROM_MEM[1192] <= 8'h85;
ROM_MEM[1193] <= 8'h04;
ROM_MEM[1194] <= 8'h10;
ROM_MEM[1195] <= 8'h26;
ROM_MEM[1196] <= 8'h00;
ROM_MEM[1197] <= 8'h9C;
ROM_MEM[1198] <= 8'hCC;
ROM_MEM[1199] <= 8'h06;
ROM_MEM[1200] <= 8'h90;
ROM_MEM[1201] <= 8'hFD;
ROM_MEM[1202] <= 8'h50;
ROM_MEM[1203] <= 8'h02;
ROM_MEM[1204] <= 8'hCC;
ROM_MEM[1205] <= 8'h05;
ROM_MEM[1206] <= 8'hA0;
ROM_MEM[1207] <= 8'hFD;
ROM_MEM[1208] <= 8'h50;
ROM_MEM[1209] <= 8'h04;
ROM_MEM[1210] <= 8'hFC;
ROM_MEM[1211] <= 8'h50;
ROM_MEM[1212] <= 8'h00;
ROM_MEM[1213] <= 8'h83;
ROM_MEM[1214] <= 8'h01;
ROM_MEM[1215] <= 8'h00;
ROM_MEM[1216] <= 8'h2A;
ROM_MEM[1217] <= 8'h03;
ROM_MEM[1218] <= 8'hCC;
ROM_MEM[1219] <= 8'h00;
ROM_MEM[1220] <= 8'h00;
ROM_MEM[1221] <= 8'hFD;
ROM_MEM[1222] <= 8'h50;
ROM_MEM[1223] <= 8'h00;
ROM_MEM[1224] <= 8'h86;
ROM_MEM[1225] <= 8'h86;
ROM_MEM[1226] <= 8'hBD;
ROM_MEM[1227] <= 8'hCD;
ROM_MEM[1228] <= 8'hBA;
ROM_MEM[1229] <= 8'hFC;
ROM_MEM[1230] <= 8'h50;
ROM_MEM[1231] <= 8'h1A;
ROM_MEM[1232] <= 8'hF3;
ROM_MEM[1233] <= 8'h50;
ROM_MEM[1234] <= 8'h02;
ROM_MEM[1235] <= 8'hC3;
ROM_MEM[1236] <= 8'h00;
ROM_MEM[1237] <= 8'h0A;
ROM_MEM[1238] <= 8'hB3;
ROM_MEM[1239] <= 8'h50;
ROM_MEM[1240] <= 8'h78;
ROM_MEM[1241] <= 8'h10;
ROM_MEM[1242] <= 8'h2D;
ROM_MEM[1243] <= 8'h00;
ROM_MEM[1244] <= 8'h6D;
ROM_MEM[1245] <= 8'h47;
ROM_MEM[1246] <= 8'h56;
ROM_MEM[1247] <= 8'h83;
ROM_MEM[1248] <= 8'h00;
ROM_MEM[1249] <= 8'h0A;
ROM_MEM[1250] <= 8'hB3;
ROM_MEM[1251] <= 8'h50;
ROM_MEM[1252] <= 8'h02;
ROM_MEM[1253] <= 8'h10;
ROM_MEM[1254] <= 8'h2E;
ROM_MEM[1255] <= 8'h00;
ROM_MEM[1256] <= 8'h61;
ROM_MEM[1257] <= 8'hFC;
ROM_MEM[1258] <= 8'h50;
ROM_MEM[1259] <= 8'h7A;
ROM_MEM[1260] <= 8'hB3;
ROM_MEM[1261] <= 8'h50;
ROM_MEM[1262] <= 8'h1C;
ROM_MEM[1263] <= 8'h2B;
ROM_MEM[1264] <= 8'h59;
ROM_MEM[1265] <= 8'hB3;
ROM_MEM[1266] <= 8'h50;
ROM_MEM[1267] <= 8'h04;
ROM_MEM[1268] <= 8'h2E;
ROM_MEM[1269] <= 8'h54;
ROM_MEM[1270] <= 8'hA6;
ROM_MEM[1271] <= 8'h04;
ROM_MEM[1272] <= 8'h81;
ROM_MEM[1273] <= 8'h03;
ROM_MEM[1274] <= 8'h26;
ROM_MEM[1275] <= 8'h0E;
ROM_MEM[1276] <= 8'hFC;
ROM_MEM[1277] <= 8'h50;
ROM_MEM[1278] <= 8'h7C;
ROM_MEM[1279] <= 8'h10;
ROM_MEM[1280] <= 8'h93;
ROM_MEM[1281] <= 8'hC8;
ROM_MEM[1282] <= 8'h24;
ROM_MEM[1283] <= 8'h04;
ROM_MEM[1284] <= 8'hDD;
ROM_MEM[1285] <= 8'hC8;
ROM_MEM[1286] <= 8'h9F;
ROM_MEM[1287] <= 8'hC6;
ROM_MEM[1288] <= 8'h20;
ROM_MEM[1289] <= 8'h40;
ROM_MEM[1290] <= 8'hCC;
ROM_MEM[1291] <= 8'h4C;
ROM_MEM[1292] <= 8'hE0;
ROM_MEM[1293] <= 8'hFD;
ROM_MEM[1294] <= 8'h50;
ROM_MEM[1295] <= 8'h02;
ROM_MEM[1296] <= 8'h86;
ROM_MEM[1297] <= 8'h86;
ROM_MEM[1298] <= 8'hBD;
ROM_MEM[1299] <= 8'hCD;
ROM_MEM[1300] <= 8'hBA;
ROM_MEM[1301] <= 8'hFC;
ROM_MEM[1302] <= 8'h50;
ROM_MEM[1303] <= 8'h7A;
ROM_MEM[1304] <= 8'hC3;
ROM_MEM[1305] <= 8'h00;
ROM_MEM[1306] <= 8'h0A;
ROM_MEM[1307] <= 8'hB3;
ROM_MEM[1308] <= 8'h50;
ROM_MEM[1309] <= 8'h1C;
ROM_MEM[1310] <= 8'hB3;
ROM_MEM[1311] <= 8'h50;
ROM_MEM[1312] <= 8'h02;
ROM_MEM[1313] <= 8'h2D;
ROM_MEM[1314] <= 8'h1B;
ROM_MEM[1315] <= 8'hCE;
ROM_MEM[1316] <= 8'h49;
ROM_MEM[1317] <= 8'hC2;
ROM_MEM[1318] <= 8'hE6;
ROM_MEM[1319] <= 8'h06;
ROM_MEM[1320] <= 8'h33;
ROM_MEM[1321] <= 8'hC5;
ROM_MEM[1322] <= 8'hA6;
ROM_MEM[1323] <= 8'hC4;
ROM_MEM[1324] <= 8'h85;
ROM_MEM[1325] <= 8'h04;
ROM_MEM[1326] <= 8'h26;
ROM_MEM[1327] <= 8'h1A;
ROM_MEM[1328] <= 8'hFC;
ROM_MEM[1329] <= 8'h50;
ROM_MEM[1330] <= 8'h7C;
ROM_MEM[1331] <= 8'h10;
ROM_MEM[1332] <= 8'h93;
ROM_MEM[1333] <= 8'hC8;
ROM_MEM[1334] <= 8'h24;
ROM_MEM[1335] <= 8'h04;
ROM_MEM[1336] <= 8'hDD;
ROM_MEM[1337] <= 8'hC8;
ROM_MEM[1338] <= 8'h9F;
ROM_MEM[1339] <= 8'hC6;
ROM_MEM[1340] <= 8'h20;
ROM_MEM[1341] <= 8'h0C;
ROM_MEM[1342] <= 8'hFC;
ROM_MEM[1343] <= 8'h50;
ROM_MEM[1344] <= 8'h7C;
ROM_MEM[1345] <= 8'h10;
ROM_MEM[1346] <= 8'h93;
ROM_MEM[1347] <= 8'hD0;
ROM_MEM[1348] <= 8'h24;
ROM_MEM[1349] <= 8'h04;
ROM_MEM[1350] <= 8'hDD;
ROM_MEM[1351] <= 8'hD0;
ROM_MEM[1352] <= 8'h9F;
ROM_MEM[1353] <= 8'hCE;
ROM_MEM[1354] <= 8'h39;
ROM_MEM[1355] <= 8'h9E;
ROM_MEM[1356] <= 8'hC6;
ROM_MEM[1357] <= 8'hEC;
ROM_MEM[1358] <= 8'h84;
ROM_MEM[1359] <= 8'hB3;
ROM_MEM[1360] <= 8'h50;
ROM_MEM[1361] <= 8'h98;
ROM_MEM[1362] <= 8'h84;
ROM_MEM[1363] <= 8'h7F;
ROM_MEM[1364] <= 8'hF3;
ROM_MEM[1365] <= 8'h50;
ROM_MEM[1366] <= 8'h98;
ROM_MEM[1367] <= 8'hFD;
ROM_MEM[1368] <= 8'h50;
ROM_MEM[1369] <= 8'h18;
ROM_MEM[1370] <= 8'hEC;
ROM_MEM[1371] <= 8'h02;
ROM_MEM[1372] <= 8'hFD;
ROM_MEM[1373] <= 8'h50;
ROM_MEM[1374] <= 8'h1A;
ROM_MEM[1375] <= 8'hCE;
ROM_MEM[1376] <= 8'h49;
ROM_MEM[1377] <= 8'hC2;
ROM_MEM[1378] <= 8'hE6;
ROM_MEM[1379] <= 8'h06;
ROM_MEM[1380] <= 8'h33;
ROM_MEM[1381] <= 8'hC5;
ROM_MEM[1382] <= 8'hA6;
ROM_MEM[1383] <= 8'hC4;
ROM_MEM[1384] <= 8'h8A;
ROM_MEM[1385] <= 8'h04;
ROM_MEM[1386] <= 8'hA7;
ROM_MEM[1387] <= 8'hC4;
ROM_MEM[1388] <= 8'hA6;
ROM_MEM[1389] <= 8'h04;
ROM_MEM[1390] <= 8'h81;
ROM_MEM[1391] <= 8'h03;
ROM_MEM[1392] <= 8'h26;
ROM_MEM[1393] <= 8'h0E;
ROM_MEM[1394] <= 8'hCC;
ROM_MEM[1395] <= 8'h02;
ROM_MEM[1396] <= 8'hD0;
ROM_MEM[1397] <= 8'hFD;
ROM_MEM[1398] <= 8'h50;
ROM_MEM[1399] <= 8'h1C;
ROM_MEM[1400] <= 8'hBD;
ROM_MEM[1401] <= 8'hB8;
ROM_MEM[1402] <= 8'h52;
ROM_MEM[1403] <= 8'hBD;
ROM_MEM[1404] <= 8'h97;
ROM_MEM[1405] <= 8'hF7;
ROM_MEM[1406] <= 8'h20;
ROM_MEM[1407] <= 8'h0C;
ROM_MEM[1408] <= 8'hCC;
ROM_MEM[1409] <= 8'h54;
ROM_MEM[1410] <= 8'h60;
ROM_MEM[1411] <= 8'hFD;
ROM_MEM[1412] <= 8'h50;
ROM_MEM[1413] <= 8'h1C;
ROM_MEM[1414] <= 8'hBD;
ROM_MEM[1415] <= 8'hB8;
ROM_MEM[1416] <= 8'h5E;
ROM_MEM[1417] <= 8'hBD;
ROM_MEM[1418] <= 8'h97;
ROM_MEM[1419] <= 8'h3A;
ROM_MEM[1420] <= 8'hBD;
ROM_MEM[1421] <= 8'hBD;
ROM_MEM[1422] <= 8'hFD;
ROM_MEM[1423] <= 8'h39;
ROM_MEM[1424] <= 8'h39;
ROM_MEM[1425] <= 8'h96;
ROM_MEM[1426] <= 8'h60;
ROM_MEM[1427] <= 8'h2D;
ROM_MEM[1428] <= 8'h1D;
ROM_MEM[1429] <= 8'h9E;
ROM_MEM[1430] <= 8'h64;
ROM_MEM[1431] <= 8'hCE;
ROM_MEM[1432] <= 8'h49;
ROM_MEM[1433] <= 8'hC2;
ROM_MEM[1434] <= 8'hE6;
ROM_MEM[1435] <= 8'h06;
ROM_MEM[1436] <= 8'h33;
ROM_MEM[1437] <= 8'hC5;
ROM_MEM[1438] <= 8'hA6;
ROM_MEM[1439] <= 8'hC4;
ROM_MEM[1440] <= 8'h85;
ROM_MEM[1441] <= 8'h04;
ROM_MEM[1442] <= 8'h26;
ROM_MEM[1443] <= 8'h0E;
ROM_MEM[1444] <= 8'hA6;
ROM_MEM[1445] <= 8'h04;
ROM_MEM[1446] <= 8'h81;
ROM_MEM[1447] <= 8'h02;
ROM_MEM[1448] <= 8'h10;
ROM_MEM[1449] <= 8'h27;
ROM_MEM[1450] <= 8'h00;
ROM_MEM[1451] <= 8'h5C;
ROM_MEM[1452] <= 8'h10;
ROM_MEM[1453] <= 8'h22;
ROM_MEM[1454] <= 8'h00;
ROM_MEM[1455] <= 8'hA5;
ROM_MEM[1456] <= 8'h20;
ROM_MEM[1457] <= 8'h01;
ROM_MEM[1458] <= 8'h39;
ROM_MEM[1459] <= 8'hCC;
ROM_MEM[1460] <= 8'h40;
ROM_MEM[1461] <= 8'h00;
ROM_MEM[1462] <= 8'hB3;
ROM_MEM[1463] <= 8'h50;
ROM_MEM[1464] <= 8'h7C;
ROM_MEM[1465] <= 8'h58;
ROM_MEM[1466] <= 8'h49;
ROM_MEM[1467] <= 8'hFD;
ROM_MEM[1468] <= 8'h50;
ROM_MEM[1469] <= 8'h00;
ROM_MEM[1470] <= 8'hCC;
ROM_MEM[1471] <= 8'h29;
ROM_MEM[1472] <= 8'h40;
ROM_MEM[1473] <= 8'hFD;
ROM_MEM[1474] <= 8'h50;
ROM_MEM[1475] <= 8'h04;
ROM_MEM[1476] <= 8'hCC;
ROM_MEM[1477] <= 8'h02;
ROM_MEM[1478] <= 8'hD0;
ROM_MEM[1479] <= 8'hFD;
ROM_MEM[1480] <= 8'h50;
ROM_MEM[1481] <= 8'h02;
ROM_MEM[1482] <= 8'h86;
ROM_MEM[1483] <= 8'h86;
ROM_MEM[1484] <= 8'hBD;
ROM_MEM[1485] <= 8'hCD;
ROM_MEM[1486] <= 8'hBA;
ROM_MEM[1487] <= 8'hFC;
ROM_MEM[1488] <= 8'h50;
ROM_MEM[1489] <= 8'h04;
ROM_MEM[1490] <= 8'hB3;
ROM_MEM[1491] <= 8'h50;
ROM_MEM[1492] <= 8'h44;
ROM_MEM[1493] <= 8'h2C;
ROM_MEM[1494] <= 8'h07;
ROM_MEM[1495] <= 8'hA6;
ROM_MEM[1496] <= 8'hC4;
ROM_MEM[1497] <= 8'h8A;
ROM_MEM[1498] <= 8'h08;
ROM_MEM[1499] <= 8'hA7;
ROM_MEM[1500] <= 8'hC4;
ROM_MEM[1501] <= 8'h39;
ROM_MEM[1502] <= 8'hB3;
ROM_MEM[1503] <= 8'h50;
ROM_MEM[1504] <= 8'h02;
ROM_MEM[1505] <= 8'h2F;
ROM_MEM[1506] <= 8'h06;
ROM_MEM[1507] <= 8'hA6;
ROM_MEM[1508] <= 8'hC4;
ROM_MEM[1509] <= 8'h85;
ROM_MEM[1510] <= 8'h08;
ROM_MEM[1511] <= 8'h27;
ROM_MEM[1512] <= 8'h1E;
ROM_MEM[1513] <= 8'hA6;
ROM_MEM[1514] <= 8'hC4;
ROM_MEM[1515] <= 8'h84;
ROM_MEM[1516] <= 8'hF7;
ROM_MEM[1517] <= 8'hA7;
ROM_MEM[1518] <= 8'hC4;
ROM_MEM[1519] <= 8'hB6;
ROM_MEM[1520] <= 8'h47;
ROM_MEM[1521] <= 8'h03;
ROM_MEM[1522] <= 8'h2A;
ROM_MEM[1523] <= 8'h03;
ROM_MEM[1524] <= 8'hBD;
ROM_MEM[1525] <= 8'hA7;
ROM_MEM[1526] <= 8'hB6;
ROM_MEM[1527] <= 8'hB6;
ROM_MEM[1528] <= 8'h47;
ROM_MEM[1529] <= 8'h03;
ROM_MEM[1530] <= 8'h2A;
ROM_MEM[1531] <= 8'h03;
ROM_MEM[1532] <= 8'hBD;
ROM_MEM[1533] <= 8'hA7;
ROM_MEM[1534] <= 8'hC8;
ROM_MEM[1535] <= 8'hB6;
ROM_MEM[1536] <= 8'h47;
ROM_MEM[1537] <= 8'h03;
ROM_MEM[1538] <= 8'h2A;
ROM_MEM[1539] <= 8'h03;
ROM_MEM[1540] <= 8'hBD;
ROM_MEM[1541] <= 8'hA7;
ROM_MEM[1542] <= 8'hBF;
ROM_MEM[1543] <= 8'h39;
ROM_MEM[1544] <= 8'hCC;
ROM_MEM[1545] <= 8'h40;
ROM_MEM[1546] <= 8'h00;
ROM_MEM[1547] <= 8'hB3;
ROM_MEM[1548] <= 8'h50;
ROM_MEM[1549] <= 8'h7C;
ROM_MEM[1550] <= 8'h58;
ROM_MEM[1551] <= 8'h49;
ROM_MEM[1552] <= 8'hFD;
ROM_MEM[1553] <= 8'h50;
ROM_MEM[1554] <= 8'h00;
ROM_MEM[1555] <= 8'hCC;
ROM_MEM[1556] <= 8'h29;
ROM_MEM[1557] <= 8'h40;
ROM_MEM[1558] <= 8'hFD;
ROM_MEM[1559] <= 8'h50;
ROM_MEM[1560] <= 8'h04;
ROM_MEM[1561] <= 8'hCC;
ROM_MEM[1562] <= 8'h02;
ROM_MEM[1563] <= 8'hD0;
ROM_MEM[1564] <= 8'hFD;
ROM_MEM[1565] <= 8'h50;
ROM_MEM[1566] <= 8'h02;
ROM_MEM[1567] <= 8'h86;
ROM_MEM[1568] <= 8'h86;
ROM_MEM[1569] <= 8'hBD;
ROM_MEM[1570] <= 8'hCD;
ROM_MEM[1571] <= 8'hBA;
ROM_MEM[1572] <= 8'hFC;
ROM_MEM[1573] <= 8'h50;
ROM_MEM[1574] <= 8'h04;
ROM_MEM[1575] <= 8'hB3;
ROM_MEM[1576] <= 8'h50;
ROM_MEM[1577] <= 8'h44;
ROM_MEM[1578] <= 8'h2C;
ROM_MEM[1579] <= 8'h07;
ROM_MEM[1580] <= 8'hA6;
ROM_MEM[1581] <= 8'hC4;
ROM_MEM[1582] <= 8'h8A;
ROM_MEM[1583] <= 8'h08;
ROM_MEM[1584] <= 8'hA7;
ROM_MEM[1585] <= 8'hC4;
ROM_MEM[1586] <= 8'h39;
ROM_MEM[1587] <= 8'hB3;
ROM_MEM[1588] <= 8'h50;
ROM_MEM[1589] <= 8'h02;
ROM_MEM[1590] <= 8'h2F;
ROM_MEM[1591] <= 8'h06;
ROM_MEM[1592] <= 8'hA6;
ROM_MEM[1593] <= 8'hC4;
ROM_MEM[1594] <= 8'h85;
ROM_MEM[1595] <= 8'h08;
ROM_MEM[1596] <= 8'h27;
ROM_MEM[1597] <= 8'h16;
ROM_MEM[1598] <= 8'hA6;
ROM_MEM[1599] <= 8'hC4;
ROM_MEM[1600] <= 8'h84;
ROM_MEM[1601] <= 8'hF7;
ROM_MEM[1602] <= 8'hA7;
ROM_MEM[1603] <= 8'hC4;
ROM_MEM[1604] <= 8'hB6;
ROM_MEM[1605] <= 8'h47;
ROM_MEM[1606] <= 8'h03;
ROM_MEM[1607] <= 8'h2A;
ROM_MEM[1608] <= 8'h03;
ROM_MEM[1609] <= 8'hBD;
ROM_MEM[1610] <= 8'hA7;
ROM_MEM[1611] <= 8'hC8;
ROM_MEM[1612] <= 8'hB6;
ROM_MEM[1613] <= 8'h47;
ROM_MEM[1614] <= 8'h03;
ROM_MEM[1615] <= 8'h2A;
ROM_MEM[1616] <= 8'h03;
ROM_MEM[1617] <= 8'hBD;
ROM_MEM[1618] <= 8'hA7;
ROM_MEM[1619] <= 8'hBF;
ROM_MEM[1620] <= 8'h39;
ROM_MEM[1621] <= 8'h86;
ROM_MEM[1622] <= 8'h40;
ROM_MEM[1623] <= 8'hB0;
ROM_MEM[1624] <= 8'h50;
ROM_MEM[1625] <= 8'h7C;
ROM_MEM[1626] <= 8'hB1;
ROM_MEM[1627] <= 8'h47;
ROM_MEM[1628] <= 8'h03;
ROM_MEM[1629] <= 8'h25;
ROM_MEM[1630] <= 8'h15;
ROM_MEM[1631] <= 8'hB6;
ROM_MEM[1632] <= 8'h47;
ROM_MEM[1633] <= 8'h03;
ROM_MEM[1634] <= 8'h81;
ROM_MEM[1635] <= 8'h50;
ROM_MEM[1636] <= 8'h24;
ROM_MEM[1637] <= 8'h03;
ROM_MEM[1638] <= 8'h7E;
ROM_MEM[1639] <= 8'hA7;
ROM_MEM[1640] <= 8'h28;
ROM_MEM[1641] <= 8'hB6;
ROM_MEM[1642] <= 8'h47;
ROM_MEM[1643] <= 8'h03;
ROM_MEM[1644] <= 8'h2A;
ROM_MEM[1645] <= 8'h03;
ROM_MEM[1646] <= 8'h7E;
ROM_MEM[1647] <= 8'hA7;
ROM_MEM[1648] <= 8'h28;
ROM_MEM[1649] <= 8'h7E;
ROM_MEM[1650] <= 8'hA7;
ROM_MEM[1651] <= 8'h28;
ROM_MEM[1652] <= 8'h39;
ROM_MEM[1653] <= 8'hA8;
ROM_MEM[1654] <= 8'h6B;
ROM_MEM[1655] <= 8'hA8;
ROM_MEM[1656] <= 8'h75;
ROM_MEM[1657] <= 8'hA8;
ROM_MEM[1658] <= 8'hA7;
ROM_MEM[1659] <= 8'hA8;
ROM_MEM[1660] <= 8'hDA;
ROM_MEM[1661] <= 8'hA8;
ROM_MEM[1662] <= 8'hE6;
ROM_MEM[1663] <= 8'hA8;
ROM_MEM[1664] <= 8'hF9;
ROM_MEM[1665] <= 8'hAA;
ROM_MEM[1666] <= 8'h00;
ROM_MEM[1667] <= 8'hA9;
ROM_MEM[1668] <= 8'h46;
ROM_MEM[1669] <= 8'hA9;
ROM_MEM[1670] <= 8'hA3;
ROM_MEM[1671] <= 8'hAA;
ROM_MEM[1672] <= 8'h86;
ROM_MEM[1673] <= 8'hAA;
ROM_MEM[1674] <= 8'hB5;
ROM_MEM[1675] <= 8'hDF;
ROM_MEM[1676] <= 8'hA8;
ROM_MEM[1677] <= 8'hC6;
ROM_MEM[1678] <= 8'h40;
ROM_MEM[1679] <= 8'hE7;
ROM_MEM[1680] <= 8'h45;
ROM_MEM[1681] <= 8'hC6;
ROM_MEM[1682] <= 8'h01;
ROM_MEM[1683] <= 8'hE7;
ROM_MEM[1684] <= 8'h43;
ROM_MEM[1685] <= 8'hC6;
ROM_MEM[1686] <= 8'h01;
ROM_MEM[1687] <= 8'hE7;
ROM_MEM[1688] <= 8'h44;
ROM_MEM[1689] <= 8'hB6;
ROM_MEM[1690] <= 8'h4B;
ROM_MEM[1691] <= 8'h3C;
ROM_MEM[1692] <= 8'h2F;
ROM_MEM[1693] <= 8'h0D;
ROM_MEM[1694] <= 8'hBC;
ROM_MEM[1695] <= 8'h4B;
ROM_MEM[1696] <= 8'h32;
ROM_MEM[1697] <= 8'h26;
ROM_MEM[1698] <= 8'h08;
ROM_MEM[1699] <= 8'h7A;
ROM_MEM[1700] <= 8'h4B;
ROM_MEM[1701] <= 8'h3C;
ROM_MEM[1702] <= 8'h26;
ROM_MEM[1703] <= 8'h03;
ROM_MEM[1704] <= 8'hBD;
ROM_MEM[1705] <= 8'hBD;
ROM_MEM[1706] <= 8'h4E;
ROM_MEM[1707] <= 8'hEE;
ROM_MEM[1708] <= 8'hC4;
ROM_MEM[1709] <= 8'hAE;
ROM_MEM[1710] <= 8'h84;
ROM_MEM[1711] <= 8'hEC;
ROM_MEM[1712] <= 8'h08;
ROM_MEM[1713] <= 8'hB3;
ROM_MEM[1714] <= 8'h50;
ROM_MEM[1715] <= 8'h98;
ROM_MEM[1716] <= 8'hED;
ROM_MEM[1717] <= 8'hC4;
ROM_MEM[1718] <= 8'hEC;
ROM_MEM[1719] <= 8'h0A;
ROM_MEM[1720] <= 8'hB3;
ROM_MEM[1721] <= 8'h50;
ROM_MEM[1722] <= 8'h9A;
ROM_MEM[1723] <= 8'hED;
ROM_MEM[1724] <= 8'h42;
ROM_MEM[1725] <= 8'hEC;
ROM_MEM[1726] <= 8'h0C;
ROM_MEM[1727] <= 8'hB3;
ROM_MEM[1728] <= 8'h50;
ROM_MEM[1729] <= 8'h9C;
ROM_MEM[1730] <= 8'hED;
ROM_MEM[1731] <= 8'h44;
ROM_MEM[1732] <= 8'hBD;
ROM_MEM[1733] <= 8'hBE;
ROM_MEM[1734] <= 8'h02;
ROM_MEM[1735] <= 8'h39;
ROM_MEM[1736] <= 8'h49;
ROM_MEM[1737] <= 8'h69;
ROM_MEM[1738] <= 8'h49;
ROM_MEM[1739] <= 8'h69;
ROM_MEM[1740] <= 8'h49;
ROM_MEM[1741] <= 8'h63;
ROM_MEM[1742] <= 8'h49;
ROM_MEM[1743] <= 8'h63;
ROM_MEM[1744] <= 8'h49;
ROM_MEM[1745] <= 8'h5D;
ROM_MEM[1746] <= 8'h49;
ROM_MEM[1747] <= 8'h5D;
ROM_MEM[1748] <= 8'h49;
ROM_MEM[1749] <= 8'h57;
ROM_MEM[1750] <= 8'h49;
ROM_MEM[1751] <= 8'h57;
ROM_MEM[1752] <= 8'h49;
ROM_MEM[1753] <= 8'h51;
ROM_MEM[1754] <= 8'h49;
ROM_MEM[1755] <= 8'h51;
ROM_MEM[1756] <= 8'h49;
ROM_MEM[1757] <= 8'h4B;
ROM_MEM[1758] <= 8'h49;
ROM_MEM[1759] <= 8'h4B;
ROM_MEM[1760] <= 8'hF6;
ROM_MEM[1761] <= 8'h4B;
ROM_MEM[1762] <= 8'h19;
ROM_MEM[1763] <= 8'hC1;
ROM_MEM[1764] <= 8'h0C;
ROM_MEM[1765] <= 8'h25;
ROM_MEM[1766] <= 8'h05;
ROM_MEM[1767] <= 8'h8E;
ROM_MEM[1768] <= 8'hA6;
ROM_MEM[1769] <= 8'hDE;
ROM_MEM[1770] <= 8'h20;
ROM_MEM[1771] <= 8'h06;
ROM_MEM[1772] <= 8'h58;
ROM_MEM[1773] <= 8'h8E;
ROM_MEM[1774] <= 8'hA6;
ROM_MEM[1775] <= 8'hC8;
ROM_MEM[1776] <= 8'hAE;
ROM_MEM[1777] <= 8'h85;
ROM_MEM[1778] <= 8'h20;
ROM_MEM[1779] <= 8'h14;
ROM_MEM[1780] <= 8'hF6;
ROM_MEM[1781] <= 8'h4B;
ROM_MEM[1782] <= 8'h19;
ROM_MEM[1783] <= 8'hC1;
ROM_MEM[1784] <= 8'h07;
ROM_MEM[1785] <= 8'h23;
ROM_MEM[1786] <= 8'h02;
ROM_MEM[1787] <= 8'hC6;
ROM_MEM[1788] <= 8'h07;
ROM_MEM[1789] <= 8'h58;
ROM_MEM[1790] <= 8'h8E;
ROM_MEM[1791] <= 8'hA7;
ROM_MEM[1792] <= 8'h18;
ROM_MEM[1793] <= 8'hAE;
ROM_MEM[1794] <= 8'h85;
ROM_MEM[1795] <= 8'h20;
ROM_MEM[1796] <= 8'h03;
ROM_MEM[1797] <= 8'h8E;
ROM_MEM[1798] <= 8'h49;
ROM_MEM[1799] <= 8'h4B;
ROM_MEM[1800] <= 8'h9F;
ROM_MEM[1801] <= 8'hA8;
ROM_MEM[1802] <= 8'hA6;
ROM_MEM[1803] <= 8'h03;
ROM_MEM[1804] <= 8'h27;
ROM_MEM[1805] <= 8'h09;
ROM_MEM[1806] <= 8'h30;
ROM_MEM[1807] <= 8'h06;
ROM_MEM[1808] <= 8'h8C;
ROM_MEM[1809] <= 8'h49;
ROM_MEM[1810] <= 8'h6F;
ROM_MEM[1811] <= 8'h25;
ROM_MEM[1812] <= 8'hF3;
ROM_MEM[1813] <= 8'h32;
ROM_MEM[1814] <= 8'h62;
ROM_MEM[1815] <= 8'h39;
ROM_MEM[1816] <= 8'h49;
ROM_MEM[1817] <= 8'h69;
ROM_MEM[1818] <= 8'h49;
ROM_MEM[1819] <= 8'h69;
ROM_MEM[1820] <= 8'h49;
ROM_MEM[1821] <= 8'h63;
ROM_MEM[1822] <= 8'h49;
ROM_MEM[1823] <= 8'h63;
ROM_MEM[1824] <= 8'h49;
ROM_MEM[1825] <= 8'h5D;
ROM_MEM[1826] <= 8'h49;
ROM_MEM[1827] <= 8'h5D;
ROM_MEM[1828] <= 8'h49;
ROM_MEM[1829] <= 8'h5D;
ROM_MEM[1830] <= 8'h49;
ROM_MEM[1831] <= 8'h57;
ROM_MEM[1832] <= 8'hBD;
ROM_MEM[1833] <= 8'hA6;
ROM_MEM[1834] <= 8'hE0;
ROM_MEM[1835] <= 8'h86;
ROM_MEM[1836] <= 8'h70;
ROM_MEM[1837] <= 8'hA7;
ROM_MEM[1838] <= 8'h05;
ROM_MEM[1839] <= 8'h86;
ROM_MEM[1840] <= 8'h05;
ROM_MEM[1841] <= 8'hA7;
ROM_MEM[1842] <= 8'h03;
ROM_MEM[1843] <= 8'hDE;
ROM_MEM[1844] <= 8'h64;
ROM_MEM[1845] <= 8'h9F;
ROM_MEM[1846] <= 8'h01;
ROM_MEM[1847] <= 8'hEC;
ROM_MEM[1848] <= 8'h42;
ROM_MEM[1849] <= 8'hB3;
ROM_MEM[1850] <= 8'h50;
ROM_MEM[1851] <= 8'h9A;
ROM_MEM[1852] <= 8'h2B;
ROM_MEM[1853] <= 8'h04;
ROM_MEM[1854] <= 8'h86;
ROM_MEM[1855] <= 8'h08;
ROM_MEM[1856] <= 8'h20;
ROM_MEM[1857] <= 8'h02;
ROM_MEM[1858] <= 8'h86;
ROM_MEM[1859] <= 8'h07;
ROM_MEM[1860] <= 8'hA7;
ROM_MEM[1861] <= 8'h04;
ROM_MEM[1862] <= 8'hAE;
ROM_MEM[1863] <= 8'h84;
ROM_MEM[1864] <= 8'hA6;
ROM_MEM[1865] <= 8'hC4;
ROM_MEM[1866] <= 8'hB0;
ROM_MEM[1867] <= 8'h50;
ROM_MEM[1868] <= 8'h98;
ROM_MEM[1869] <= 8'h84;
ROM_MEM[1870] <= 8'h80;
ROM_MEM[1871] <= 8'hA8;
ROM_MEM[1872] <= 8'hC4;
ROM_MEM[1873] <= 8'hE6;
ROM_MEM[1874] <= 8'h41;
ROM_MEM[1875] <= 8'hED;
ROM_MEM[1876] <= 8'h84;
ROM_MEM[1877] <= 8'hEC;
ROM_MEM[1878] <= 8'h42;
ROM_MEM[1879] <= 8'hED;
ROM_MEM[1880] <= 8'h02;
ROM_MEM[1881] <= 8'hCC;
ROM_MEM[1882] <= 8'h02;
ROM_MEM[1883] <= 8'h00;
ROM_MEM[1884] <= 8'hED;
ROM_MEM[1885] <= 8'h04;
ROM_MEM[1886] <= 8'hEC;
ROM_MEM[1887] <= 8'h02;
ROM_MEM[1888] <= 8'hB3;
ROM_MEM[1889] <= 8'h50;
ROM_MEM[1890] <= 8'h9A;
ROM_MEM[1891] <= 8'hA7;
ROM_MEM[1892] <= 8'h06;
ROM_MEM[1893] <= 8'h2A;
ROM_MEM[1894] <= 8'h04;
ROM_MEM[1895] <= 8'h43;
ROM_MEM[1896] <= 8'h50;
ROM_MEM[1897] <= 8'h82;
ROM_MEM[1898] <= 8'hFF;
ROM_MEM[1899] <= 8'hFD;
ROM_MEM[1900] <= 8'h47;
ROM_MEM[1901] <= 8'h06;
ROM_MEM[1902] <= 8'hEC;
ROM_MEM[1903] <= 8'h84;
ROM_MEM[1904] <= 8'hB3;
ROM_MEM[1905] <= 8'h50;
ROM_MEM[1906] <= 8'h98;
ROM_MEM[1907] <= 8'hFD;
ROM_MEM[1908] <= 8'h47;
ROM_MEM[1909] <= 8'h04;
ROM_MEM[1910] <= 8'hCC;
ROM_MEM[1911] <= 8'h02;
ROM_MEM[1912] <= 8'h00;
ROM_MEM[1913] <= 8'hFD;
ROM_MEM[1914] <= 8'h47;
ROM_MEM[1915] <= 8'h06;
ROM_MEM[1916] <= 8'hB6;
ROM_MEM[1917] <= 8'h47;
ROM_MEM[1918] <= 8'h00;
ROM_MEM[1919] <= 8'h48;
ROM_MEM[1920] <= 8'h48;
ROM_MEM[1921] <= 8'h24;
ROM_MEM[1922] <= 8'h01;
ROM_MEM[1923] <= 8'h4F;
ROM_MEM[1924] <= 8'hA7;
ROM_MEM[1925] <= 8'h07;
ROM_MEM[1926] <= 8'h96;
ROM_MEM[1927] <= 8'h7D;
ROM_MEM[1928] <= 8'hA8;
ROM_MEM[1929] <= 8'h06;
ROM_MEM[1930] <= 8'h2A;
ROM_MEM[1931] <= 8'h04;
ROM_MEM[1932] <= 8'h6F;
ROM_MEM[1933] <= 8'h06;
ROM_MEM[1934] <= 8'h20;
ROM_MEM[1935] <= 8'h22;
ROM_MEM[1936] <= 8'h96;
ROM_MEM[1937] <= 8'h7D;
ROM_MEM[1938] <= 8'h2A;
ROM_MEM[1939] <= 8'h01;
ROM_MEM[1940] <= 8'h40;
ROM_MEM[1941] <= 8'h48;
ROM_MEM[1942] <= 8'hA1;
ROM_MEM[1943] <= 8'h07;
ROM_MEM[1944] <= 8'h22;
ROM_MEM[1945] <= 8'h04;
ROM_MEM[1946] <= 8'h6F;
ROM_MEM[1947] <= 8'h06;
ROM_MEM[1948] <= 8'h20;
ROM_MEM[1949] <= 8'h14;
ROM_MEM[1950] <= 8'h86;
ROM_MEM[1951] <= 8'hFF;
ROM_MEM[1952] <= 8'hA7;
ROM_MEM[1953] <= 8'h06;
ROM_MEM[1954] <= 8'h9E;
ROM_MEM[1955] <= 8'h01;
ROM_MEM[1956] <= 8'hA6;
ROM_MEM[1957] <= 8'h04;
ROM_MEM[1958] <= 8'h81;
ROM_MEM[1959] <= 8'h08;
ROM_MEM[1960] <= 8'h26;
ROM_MEM[1961] <= 8'h04;
ROM_MEM[1962] <= 8'h86;
ROM_MEM[1963] <= 8'h07;
ROM_MEM[1964] <= 8'h20;
ROM_MEM[1965] <= 8'h02;
ROM_MEM[1966] <= 8'h86;
ROM_MEM[1967] <= 8'h08;
ROM_MEM[1968] <= 8'hA7;
ROM_MEM[1969] <= 8'h04;
ROM_MEM[1970] <= 8'hBD;
ROM_MEM[1971] <= 8'hBE;
ROM_MEM[1972] <= 8'h11;
ROM_MEM[1973] <= 8'h39;
ROM_MEM[1974] <= 8'hBD;
ROM_MEM[1975] <= 8'hA7;
ROM_MEM[1976] <= 8'h05;
ROM_MEM[1977] <= 8'h86;
ROM_MEM[1978] <= 8'h03;
ROM_MEM[1979] <= 8'hA7;
ROM_MEM[1980] <= 8'h04;
ROM_MEM[1981] <= 8'h20;
ROM_MEM[1982] <= 8'h12;
ROM_MEM[1983] <= 8'hBD;
ROM_MEM[1984] <= 8'hA7;
ROM_MEM[1985] <= 8'h05;
ROM_MEM[1986] <= 8'h86;
ROM_MEM[1987] <= 8'h04;
ROM_MEM[1988] <= 8'hA7;
ROM_MEM[1989] <= 8'h04;
ROM_MEM[1990] <= 8'h20;
ROM_MEM[1991] <= 8'h09;
ROM_MEM[1992] <= 8'hBD;
ROM_MEM[1993] <= 8'hA7;
ROM_MEM[1994] <= 8'h05;
ROM_MEM[1995] <= 8'h86;
ROM_MEM[1996] <= 8'h05;
ROM_MEM[1997] <= 8'hA7;
ROM_MEM[1998] <= 8'h04;
ROM_MEM[1999] <= 8'h20;
ROM_MEM[2000] <= 8'h00;
ROM_MEM[2001] <= 8'h86;
ROM_MEM[2002] <= 8'h70;
ROM_MEM[2003] <= 8'hA7;
ROM_MEM[2004] <= 8'h05;
ROM_MEM[2005] <= 8'h86;
ROM_MEM[2006] <= 8'h05;
ROM_MEM[2007] <= 8'hA7;
ROM_MEM[2008] <= 8'h03;
ROM_MEM[2009] <= 8'hDE;
ROM_MEM[2010] <= 8'h64;
ROM_MEM[2011] <= 8'hAE;
ROM_MEM[2012] <= 8'h84;
ROM_MEM[2013] <= 8'hA6;
ROM_MEM[2014] <= 8'hC4;
ROM_MEM[2015] <= 8'hB0;
ROM_MEM[2016] <= 8'h50;
ROM_MEM[2017] <= 8'h98;
ROM_MEM[2018] <= 8'h84;
ROM_MEM[2019] <= 8'h80;
ROM_MEM[2020] <= 8'hA8;
ROM_MEM[2021] <= 8'hC4;
ROM_MEM[2022] <= 8'hE6;
ROM_MEM[2023] <= 8'h41;
ROM_MEM[2024] <= 8'hED;
ROM_MEM[2025] <= 8'h84;
ROM_MEM[2026] <= 8'hEC;
ROM_MEM[2027] <= 8'h42;
ROM_MEM[2028] <= 8'hED;
ROM_MEM[2029] <= 8'h02;
ROM_MEM[2030] <= 8'hFC;
ROM_MEM[2031] <= 8'h50;
ROM_MEM[2032] <= 8'h44;
ROM_MEM[2033] <= 8'hED;
ROM_MEM[2034] <= 8'h04;
ROM_MEM[2035] <= 8'hBD;
ROM_MEM[2036] <= 8'hBE;
ROM_MEM[2037] <= 8'h11;
ROM_MEM[2038] <= 8'h39;
ROM_MEM[2039] <= 8'h96;
ROM_MEM[2040] <= 8'h95;
ROM_MEM[2041] <= 8'h27;
ROM_MEM[2042] <= 8'h05;
ROM_MEM[2043] <= 8'hBD;
ROM_MEM[2044] <= 8'hA7;
ROM_MEM[2045] <= 8'h05;
ROM_MEM[2046] <= 8'h20;
ROM_MEM[2047] <= 8'h03;
ROM_MEM[2048] <= 8'hBD;
ROM_MEM[2049] <= 8'hA6;
ROM_MEM[2050] <= 8'hF4;
ROM_MEM[2051] <= 8'h86;
ROM_MEM[2052] <= 8'h09;
ROM_MEM[2053] <= 8'hA7;
ROM_MEM[2054] <= 8'h04;
ROM_MEM[2055] <= 8'hEE;
ROM_MEM[2056] <= 8'h84;
ROM_MEM[2057] <= 8'h20;
ROM_MEM[2058] <= 8'h14;
ROM_MEM[2059] <= 8'h96;
ROM_MEM[2060] <= 8'h95;
ROM_MEM[2061] <= 8'h27;
ROM_MEM[2062] <= 8'h05;
ROM_MEM[2063] <= 8'hBD;
ROM_MEM[2064] <= 8'hA7;
ROM_MEM[2065] <= 8'h05;
ROM_MEM[2066] <= 8'h20;
ROM_MEM[2067] <= 8'h03;
ROM_MEM[2068] <= 8'hBD;
ROM_MEM[2069] <= 8'hA6;
ROM_MEM[2070] <= 8'hF4;
ROM_MEM[2071] <= 8'h86;
ROM_MEM[2072] <= 8'h0A;
ROM_MEM[2073] <= 8'hA7;
ROM_MEM[2074] <= 8'h04;
ROM_MEM[2075] <= 8'hEE;
ROM_MEM[2076] <= 8'h84;
ROM_MEM[2077] <= 8'h20;
ROM_MEM[2078] <= 8'h00;
ROM_MEM[2079] <= 8'hFC;
ROM_MEM[2080] <= 8'h50;
ROM_MEM[2081] <= 8'h78;
ROM_MEM[2082] <= 8'hED;
ROM_MEM[2083] <= 8'hC4;
ROM_MEM[2084] <= 8'hFC;
ROM_MEM[2085] <= 8'h50;
ROM_MEM[2086] <= 8'h7A;
ROM_MEM[2087] <= 8'hED;
ROM_MEM[2088] <= 8'h42;
ROM_MEM[2089] <= 8'hFC;
ROM_MEM[2090] <= 8'h50;
ROM_MEM[2091] <= 8'h7C;
ROM_MEM[2092] <= 8'hED;
ROM_MEM[2093] <= 8'h44;
ROM_MEM[2094] <= 8'h86;
ROM_MEM[2095] <= 8'h40;
ROM_MEM[2096] <= 8'hA7;
ROM_MEM[2097] <= 8'h05;
ROM_MEM[2098] <= 8'h86;
ROM_MEM[2099] <= 8'h05;
ROM_MEM[2100] <= 8'hA7;
ROM_MEM[2101] <= 8'h03;
ROM_MEM[2102] <= 8'hB6;
ROM_MEM[2103] <= 8'h47;
ROM_MEM[2104] <= 8'h03;
ROM_MEM[2105] <= 8'h44;
ROM_MEM[2106] <= 8'hF6;
ROM_MEM[2107] <= 8'h50;
ROM_MEM[2108] <= 8'h7C;
ROM_MEM[2109] <= 8'hC1;
ROM_MEM[2110] <= 8'hFC;
ROM_MEM[2111] <= 8'h2D;
ROM_MEM[2112] <= 8'h02;
ROM_MEM[2113] <= 8'h86;
ROM_MEM[2114] <= 8'h00;
ROM_MEM[2115] <= 8'hA7;
ROM_MEM[2116] <= 8'h46;
ROM_MEM[2117] <= 8'hBD;
ROM_MEM[2118] <= 8'hBE;
ROM_MEM[2119] <= 8'h11;
ROM_MEM[2120] <= 8'h39;
ROM_MEM[2121] <= 8'h8E;
ROM_MEM[2122] <= 8'h49;
ROM_MEM[2123] <= 8'h4B;
ROM_MEM[2124] <= 8'h9F;
ROM_MEM[2125] <= 8'hA8;
ROM_MEM[2126] <= 8'hA6;
ROM_MEM[2127] <= 8'h03;
ROM_MEM[2128] <= 8'h27;
ROM_MEM[2129] <= 8'h0F;
ROM_MEM[2130] <= 8'hE6;
ROM_MEM[2131] <= 8'h04;
ROM_MEM[2132] <= 8'h58;
ROM_MEM[2133] <= 8'hC1;
ROM_MEM[2134] <= 8'h16;
ROM_MEM[2135] <= 8'h24;
ROM_MEM[2136] <= 8'h07;
ROM_MEM[2137] <= 8'hCE;
ROM_MEM[2138] <= 8'hA6;
ROM_MEM[2139] <= 8'h75;
ROM_MEM[2140] <= 8'hAD;
ROM_MEM[2141] <= 8'hD5;
ROM_MEM[2142] <= 8'h20;
ROM_MEM[2143] <= 8'h01;
ROM_MEM[2144] <= 8'h3F;
ROM_MEM[2145] <= 8'h9E;
ROM_MEM[2146] <= 8'hA8;
ROM_MEM[2147] <= 8'h30;
ROM_MEM[2148] <= 8'h06;
ROM_MEM[2149] <= 8'h8C;
ROM_MEM[2150] <= 8'h49;
ROM_MEM[2151] <= 8'h6F;
ROM_MEM[2152] <= 8'h25;
ROM_MEM[2153] <= 8'hE2;
ROM_MEM[2154] <= 8'h39;
ROM_MEM[2155] <= 8'h6A;
ROM_MEM[2156] <= 8'h05;
ROM_MEM[2157] <= 8'h2E;
ROM_MEM[2158] <= 8'h05;
ROM_MEM[2159] <= 8'h5F;
ROM_MEM[2160] <= 8'hE7;
ROM_MEM[2161] <= 8'h03;
ROM_MEM[2162] <= 8'hE7;
ROM_MEM[2163] <= 8'h05;
ROM_MEM[2164] <= 8'h39;
ROM_MEM[2165] <= 8'h6A;
ROM_MEM[2166] <= 8'h05;
ROM_MEM[2167] <= 8'h2E;
ROM_MEM[2168] <= 8'h07;
ROM_MEM[2169] <= 8'h5F;
ROM_MEM[2170] <= 8'hE7;
ROM_MEM[2171] <= 8'h03;
ROM_MEM[2172] <= 8'hE7;
ROM_MEM[2173] <= 8'h05;
ROM_MEM[2174] <= 8'h20;
ROM_MEM[2175] <= 8'h26;
ROM_MEM[2176] <= 8'hEE;
ROM_MEM[2177] <= 8'h84;
ROM_MEM[2178] <= 8'hCC;
ROM_MEM[2179] <= 8'h00;
ROM_MEM[2180] <= 8'h00;
ROM_MEM[2181] <= 8'hA3;
ROM_MEM[2182] <= 8'hC4;
ROM_MEM[2183] <= 8'hBD;
ROM_MEM[2184] <= 8'hCD;
ROM_MEM[2185] <= 8'hA2;
ROM_MEM[2186] <= 8'hE3;
ROM_MEM[2187] <= 8'hC4;
ROM_MEM[2188] <= 8'hED;
ROM_MEM[2189] <= 8'hC4;
ROM_MEM[2190] <= 8'hCC;
ROM_MEM[2191] <= 8'h00;
ROM_MEM[2192] <= 8'h00;
ROM_MEM[2193] <= 8'hA3;
ROM_MEM[2194] <= 8'h42;
ROM_MEM[2195] <= 8'hBD;
ROM_MEM[2196] <= 8'hCD;
ROM_MEM[2197] <= 8'hA2;
ROM_MEM[2198] <= 8'hE3;
ROM_MEM[2199] <= 8'h42;
ROM_MEM[2200] <= 8'hED;
ROM_MEM[2201] <= 8'h42;
ROM_MEM[2202] <= 8'hCC;
ROM_MEM[2203] <= 8'h00;
ROM_MEM[2204] <= 8'h00;
ROM_MEM[2205] <= 8'hA3;
ROM_MEM[2206] <= 8'h44;
ROM_MEM[2207] <= 8'hBD;
ROM_MEM[2208] <= 8'hCD;
ROM_MEM[2209] <= 8'hA2;
ROM_MEM[2210] <= 8'hE3;
ROM_MEM[2211] <= 8'h44;
ROM_MEM[2212] <= 8'hED;
ROM_MEM[2213] <= 8'h44;
ROM_MEM[2214] <= 8'h39;
ROM_MEM[2215] <= 8'h6A;
ROM_MEM[2216] <= 8'h05;
ROM_MEM[2217] <= 8'h2E;
ROM_MEM[2218] <= 8'h07;
ROM_MEM[2219] <= 8'h5F;
ROM_MEM[2220] <= 8'hE7;
ROM_MEM[2221] <= 8'h03;
ROM_MEM[2222] <= 8'hE7;
ROM_MEM[2223] <= 8'h05;
ROM_MEM[2224] <= 8'h20;
ROM_MEM[2225] <= 8'h23;
ROM_MEM[2226] <= 8'hEE;
ROM_MEM[2227] <= 8'h84;
ROM_MEM[2228] <= 8'hEC;
ROM_MEM[2229] <= 8'hC4;
ROM_MEM[2230] <= 8'hBD;
ROM_MEM[2231] <= 8'hCD;
ROM_MEM[2232] <= 8'hA2;
ROM_MEM[2233] <= 8'hE3;
ROM_MEM[2234] <= 8'hC4;
ROM_MEM[2235] <= 8'h29;
ROM_MEM[2236] <= 8'h19;
ROM_MEM[2237] <= 8'hED;
ROM_MEM[2238] <= 8'hC4;
ROM_MEM[2239] <= 8'hEC;
ROM_MEM[2240] <= 8'h42;
ROM_MEM[2241] <= 8'hBD;
ROM_MEM[2242] <= 8'hCD;
ROM_MEM[2243] <= 8'hA2;
ROM_MEM[2244] <= 8'hE3;
ROM_MEM[2245] <= 8'h42;
ROM_MEM[2246] <= 8'h29;
ROM_MEM[2247] <= 8'h0E;
ROM_MEM[2248] <= 8'hED;
ROM_MEM[2249] <= 8'h42;
ROM_MEM[2250] <= 8'hEC;
ROM_MEM[2251] <= 8'h44;
ROM_MEM[2252] <= 8'hBD;
ROM_MEM[2253] <= 8'hCD;
ROM_MEM[2254] <= 8'hA2;
ROM_MEM[2255] <= 8'hE3;
ROM_MEM[2256] <= 8'h44;
ROM_MEM[2257] <= 8'h29;
ROM_MEM[2258] <= 8'h03;
ROM_MEM[2259] <= 8'hED;
ROM_MEM[2260] <= 8'h44;
ROM_MEM[2261] <= 8'h39;
ROM_MEM[2262] <= 8'h5F;
ROM_MEM[2263] <= 8'hE7;
ROM_MEM[2264] <= 8'h03;
ROM_MEM[2265] <= 8'h39;
ROM_MEM[2266] <= 8'hEE;
ROM_MEM[2267] <= 8'h84;
ROM_MEM[2268] <= 8'hCC;
ROM_MEM[2269] <= 8'hFF;
ROM_MEM[2270] <= 8'h00;
ROM_MEM[2271] <= 8'hE3;
ROM_MEM[2272] <= 8'hC4;
ROM_MEM[2273] <= 8'hED;
ROM_MEM[2274] <= 8'hC4;
ROM_MEM[2275] <= 8'h7E;
ROM_MEM[2276] <= 8'hAA;
ROM_MEM[2277] <= 8'h7D;
ROM_MEM[2278] <= 8'hEE;
ROM_MEM[2279] <= 8'h84;
ROM_MEM[2280] <= 8'hCC;
ROM_MEM[2281] <= 8'hFF;
ROM_MEM[2282] <= 8'h00;
ROM_MEM[2283] <= 8'hE3;
ROM_MEM[2284] <= 8'hC4;
ROM_MEM[2285] <= 8'hED;
ROM_MEM[2286] <= 8'hC4;
ROM_MEM[2287] <= 8'hCC;
ROM_MEM[2288] <= 8'hFF;
ROM_MEM[2289] <= 8'h00;
ROM_MEM[2290] <= 8'hE3;
ROM_MEM[2291] <= 8'h42;
ROM_MEM[2292] <= 8'hED;
ROM_MEM[2293] <= 8'h42;
ROM_MEM[2294] <= 8'h7E;
ROM_MEM[2295] <= 8'hAA;
ROM_MEM[2296] <= 8'h7D;
ROM_MEM[2297] <= 8'hEE;
ROM_MEM[2298] <= 8'h84;
ROM_MEM[2299] <= 8'hCC;
ROM_MEM[2300] <= 8'hFF;
ROM_MEM[2301] <= 8'h00;
ROM_MEM[2302] <= 8'hE3;
ROM_MEM[2303] <= 8'hC4;
ROM_MEM[2304] <= 8'hED;
ROM_MEM[2305] <= 8'hC4;
ROM_MEM[2306] <= 8'hCC;
ROM_MEM[2307] <= 8'h01;
ROM_MEM[2308] <= 8'h00;
ROM_MEM[2309] <= 8'hE3;
ROM_MEM[2310] <= 8'h42;
ROM_MEM[2311] <= 8'hED;
ROM_MEM[2312] <= 8'h42;
ROM_MEM[2313] <= 8'h7E;
ROM_MEM[2314] <= 8'hAA;
ROM_MEM[2315] <= 8'h7D;
ROM_MEM[2316] <= 8'hE6;
ROM_MEM[2317] <= 8'hC4;
ROM_MEM[2318] <= 8'hF0;
ROM_MEM[2319] <= 8'h50;
ROM_MEM[2320] <= 8'h98;
ROM_MEM[2321] <= 8'h2B;
ROM_MEM[2322] <= 8'h0C;
ROM_MEM[2323] <= 8'h4F;
ROM_MEM[2324] <= 8'hBD;
ROM_MEM[2325] <= 8'hCD;
ROM_MEM[2326] <= 8'hB5;
ROM_MEM[2327] <= 8'h43;
ROM_MEM[2328] <= 8'h50;
ROM_MEM[2329] <= 8'h82;
ROM_MEM[2330] <= 8'hFF;
ROM_MEM[2331] <= 8'hE3;
ROM_MEM[2332] <= 8'hC4;
ROM_MEM[2333] <= 8'hED;
ROM_MEM[2334] <= 8'hC4;
ROM_MEM[2335] <= 8'h39;
ROM_MEM[2336] <= 8'hCC;
ROM_MEM[2337] <= 8'h00;
ROM_MEM[2338] <= 8'h00;
ROM_MEM[2339] <= 8'hB3;
ROM_MEM[2340] <= 8'h50;
ROM_MEM[2341] <= 8'h8E;
ROM_MEM[2342] <= 8'hBD;
ROM_MEM[2343] <= 8'hCD;
ROM_MEM[2344] <= 8'hA2;
ROM_MEM[2345] <= 8'hF3;
ROM_MEM[2346] <= 8'h50;
ROM_MEM[2347] <= 8'h8E;
ROM_MEM[2348] <= 8'h2A;
ROM_MEM[2349] <= 8'h04;
ROM_MEM[2350] <= 8'hE3;
ROM_MEM[2351] <= 8'h42;
ROM_MEM[2352] <= 8'hED;
ROM_MEM[2353] <= 8'h42;
ROM_MEM[2354] <= 8'h39;
ROM_MEM[2355] <= 8'hCC;
ROM_MEM[2356] <= 8'h00;
ROM_MEM[2357] <= 8'h00;
ROM_MEM[2358] <= 8'hB3;
ROM_MEM[2359] <= 8'h50;
ROM_MEM[2360] <= 8'h8E;
ROM_MEM[2361] <= 8'hBD;
ROM_MEM[2362] <= 8'hCD;
ROM_MEM[2363] <= 8'hA2;
ROM_MEM[2364] <= 8'hF3;
ROM_MEM[2365] <= 8'h50;
ROM_MEM[2366] <= 8'h8E;
ROM_MEM[2367] <= 8'h2B;
ROM_MEM[2368] <= 8'h04;
ROM_MEM[2369] <= 8'hE3;
ROM_MEM[2370] <= 8'h42;
ROM_MEM[2371] <= 8'hED;
ROM_MEM[2372] <= 8'h42;
ROM_MEM[2373] <= 8'h39;
ROM_MEM[2374] <= 8'hEE;
ROM_MEM[2375] <= 8'h84;
ROM_MEM[2376] <= 8'hBD;
ROM_MEM[2377] <= 8'hA9;
ROM_MEM[2378] <= 8'h33;
ROM_MEM[2379] <= 8'hBD;
ROM_MEM[2380] <= 8'hA9;
ROM_MEM[2381] <= 8'h0C;
ROM_MEM[2382] <= 8'hEC;
ROM_MEM[2383] <= 8'hC4;
ROM_MEM[2384] <= 8'hB3;
ROM_MEM[2385] <= 8'h50;
ROM_MEM[2386] <= 8'h98;
ROM_MEM[2387] <= 8'hE6;
ROM_MEM[2388] <= 8'h47;
ROM_MEM[2389] <= 8'h3D;
ROM_MEM[2390] <= 8'h6D;
ROM_MEM[2391] <= 8'h46;
ROM_MEM[2392] <= 8'h26;
ROM_MEM[2393] <= 8'h04;
ROM_MEM[2394] <= 8'h43;
ROM_MEM[2395] <= 8'h50;
ROM_MEM[2396] <= 8'h82;
ROM_MEM[2397] <= 8'hFF;
ROM_MEM[2398] <= 8'hF3;
ROM_MEM[2399] <= 8'h50;
ROM_MEM[2400] <= 8'h9A;
ROM_MEM[2401] <= 8'hA3;
ROM_MEM[2402] <= 8'h42;
ROM_MEM[2403] <= 8'hC3;
ROM_MEM[2404] <= 8'h01;
ROM_MEM[2405] <= 8'h00;
ROM_MEM[2406] <= 8'h2B;
ROM_MEM[2407] <= 8'h10;
ROM_MEM[2408] <= 8'hBD;
ROM_MEM[2409] <= 8'hCD;
ROM_MEM[2410] <= 8'hA2;
ROM_MEM[2411] <= 8'h10;
ROM_MEM[2412] <= 8'h83;
ROM_MEM[2413] <= 8'h01;
ROM_MEM[2414] <= 8'h80;
ROM_MEM[2415] <= 8'h2F;
ROM_MEM[2416] <= 8'h03;
ROM_MEM[2417] <= 8'hCC;
ROM_MEM[2418] <= 8'h01;
ROM_MEM[2419] <= 8'h80;
ROM_MEM[2420] <= 8'hE3;
ROM_MEM[2421] <= 8'h42;
ROM_MEM[2422] <= 8'h20;
ROM_MEM[2423] <= 8'h0E;
ROM_MEM[2424] <= 8'hBD;
ROM_MEM[2425] <= 8'hCD;
ROM_MEM[2426] <= 8'h9E;
ROM_MEM[2427] <= 8'h10;
ROM_MEM[2428] <= 8'h83;
ROM_MEM[2429] <= 8'hFE;
ROM_MEM[2430] <= 8'h80;
ROM_MEM[2431] <= 8'h2C;
ROM_MEM[2432] <= 8'h03;
ROM_MEM[2433] <= 8'hCC;
ROM_MEM[2434] <= 8'hFE;
ROM_MEM[2435] <= 8'h80;
ROM_MEM[2436] <= 8'hE3;
ROM_MEM[2437] <= 8'h42;
ROM_MEM[2438] <= 8'hED;
ROM_MEM[2439] <= 8'h42;
ROM_MEM[2440] <= 8'hFC;
ROM_MEM[2441] <= 8'h50;
ROM_MEM[2442] <= 8'h9C;
ROM_MEM[2443] <= 8'hC3;
ROM_MEM[2444] <= 8'h01;
ROM_MEM[2445] <= 8'h00;
ROM_MEM[2446] <= 8'hA3;
ROM_MEM[2447] <= 8'h44;
ROM_MEM[2448] <= 8'h2B;
ROM_MEM[2449] <= 8'h10;
ROM_MEM[2450] <= 8'hBD;
ROM_MEM[2451] <= 8'hCD;
ROM_MEM[2452] <= 8'hA2;
ROM_MEM[2453] <= 8'h10;
ROM_MEM[2454] <= 8'h83;
ROM_MEM[2455] <= 8'h02;
ROM_MEM[2456] <= 8'h00;
ROM_MEM[2457] <= 8'h2F;
ROM_MEM[2458] <= 8'h03;
ROM_MEM[2459] <= 8'hCC;
ROM_MEM[2460] <= 8'h02;
ROM_MEM[2461] <= 8'h00;
ROM_MEM[2462] <= 8'hE3;
ROM_MEM[2463] <= 8'h44;
ROM_MEM[2464] <= 8'hED;
ROM_MEM[2465] <= 8'h44;
ROM_MEM[2466] <= 8'h39;
ROM_MEM[2467] <= 8'hEE;
ROM_MEM[2468] <= 8'h84;
ROM_MEM[2469] <= 8'hBD;
ROM_MEM[2470] <= 8'hA9;
ROM_MEM[2471] <= 8'h20;
ROM_MEM[2472] <= 8'hBD;
ROM_MEM[2473] <= 8'hA9;
ROM_MEM[2474] <= 8'h0C;
ROM_MEM[2475] <= 8'hEC;
ROM_MEM[2476] <= 8'hC4;
ROM_MEM[2477] <= 8'hB3;
ROM_MEM[2478] <= 8'h50;
ROM_MEM[2479] <= 8'h98;
ROM_MEM[2480] <= 8'hE6;
ROM_MEM[2481] <= 8'h47;
ROM_MEM[2482] <= 8'h3D;
ROM_MEM[2483] <= 8'h6D;
ROM_MEM[2484] <= 8'h46;
ROM_MEM[2485] <= 8'h27;
ROM_MEM[2486] <= 8'h04;
ROM_MEM[2487] <= 8'h43;
ROM_MEM[2488] <= 8'h50;
ROM_MEM[2489] <= 8'h82;
ROM_MEM[2490] <= 8'hFF;
ROM_MEM[2491] <= 8'hF3;
ROM_MEM[2492] <= 8'h50;
ROM_MEM[2493] <= 8'h9A;
ROM_MEM[2494] <= 8'hC3;
ROM_MEM[2495] <= 8'hFF;
ROM_MEM[2496] <= 8'h00;
ROM_MEM[2497] <= 8'hA3;
ROM_MEM[2498] <= 8'h42;
ROM_MEM[2499] <= 8'h2B;
ROM_MEM[2500] <= 8'h10;
ROM_MEM[2501] <= 8'hBD;
ROM_MEM[2502] <= 8'hCD;
ROM_MEM[2503] <= 8'h9E;
ROM_MEM[2504] <= 8'h10;
ROM_MEM[2505] <= 8'h83;
ROM_MEM[2506] <= 8'h01;
ROM_MEM[2507] <= 8'h80;
ROM_MEM[2508] <= 8'h2F;
ROM_MEM[2509] <= 8'h03;
ROM_MEM[2510] <= 8'hCC;
ROM_MEM[2511] <= 8'h01;
ROM_MEM[2512] <= 8'h80;
ROM_MEM[2513] <= 8'hE3;
ROM_MEM[2514] <= 8'h42;
ROM_MEM[2515] <= 8'h20;
ROM_MEM[2516] <= 8'h0E;
ROM_MEM[2517] <= 8'hBD;
ROM_MEM[2518] <= 8'hCD;
ROM_MEM[2519] <= 8'hA2;
ROM_MEM[2520] <= 8'h10;
ROM_MEM[2521] <= 8'h83;
ROM_MEM[2522] <= 8'hFE;
ROM_MEM[2523] <= 8'h80;
ROM_MEM[2524] <= 8'h2C;
ROM_MEM[2525] <= 8'h03;
ROM_MEM[2526] <= 8'hCC;
ROM_MEM[2527] <= 8'hFE;
ROM_MEM[2528] <= 8'h80;
ROM_MEM[2529] <= 8'hE3;
ROM_MEM[2530] <= 8'h42;
ROM_MEM[2531] <= 8'hED;
ROM_MEM[2532] <= 8'h42;
ROM_MEM[2533] <= 8'hFC;
ROM_MEM[2534] <= 8'h50;
ROM_MEM[2535] <= 8'h9C;
ROM_MEM[2536] <= 8'hC3;
ROM_MEM[2537] <= 8'h01;
ROM_MEM[2538] <= 8'h00;
ROM_MEM[2539] <= 8'hA3;
ROM_MEM[2540] <= 8'h44;
ROM_MEM[2541] <= 8'h2B;
ROM_MEM[2542] <= 8'h10;
ROM_MEM[2543] <= 8'hBD;
ROM_MEM[2544] <= 8'hCD;
ROM_MEM[2545] <= 8'hA2;
ROM_MEM[2546] <= 8'h10;
ROM_MEM[2547] <= 8'h83;
ROM_MEM[2548] <= 8'h02;
ROM_MEM[2549] <= 8'h00;
ROM_MEM[2550] <= 8'h2F;
ROM_MEM[2551] <= 8'h03;
ROM_MEM[2552] <= 8'hCC;
ROM_MEM[2553] <= 8'h02;
ROM_MEM[2554] <= 8'h00;
ROM_MEM[2555] <= 8'hE3;
ROM_MEM[2556] <= 8'h44;
ROM_MEM[2557] <= 8'hED;
ROM_MEM[2558] <= 8'h44;
ROM_MEM[2559] <= 8'h39;
ROM_MEM[2560] <= 8'hEE;
ROM_MEM[2561] <= 8'h84;
ROM_MEM[2562] <= 8'hCC;
ROM_MEM[2563] <= 8'hFF;
ROM_MEM[2564] <= 8'h00;
ROM_MEM[2565] <= 8'hE3;
ROM_MEM[2566] <= 8'hC4;
ROM_MEM[2567] <= 8'hED;
ROM_MEM[2568] <= 8'hC4;
ROM_MEM[2569] <= 8'hFC;
ROM_MEM[2570] <= 8'h50;
ROM_MEM[2571] <= 8'h9C;
ROM_MEM[2572] <= 8'hC3;
ROM_MEM[2573] <= 8'h00;
ROM_MEM[2574] <= 8'h80;
ROM_MEM[2575] <= 8'hA3;
ROM_MEM[2576] <= 8'h44;
ROM_MEM[2577] <= 8'h2B;
ROM_MEM[2578] <= 8'h10;
ROM_MEM[2579] <= 8'hBD;
ROM_MEM[2580] <= 8'hCD;
ROM_MEM[2581] <= 8'hA2;
ROM_MEM[2582] <= 8'h10;
ROM_MEM[2583] <= 8'h83;
ROM_MEM[2584] <= 8'h01;
ROM_MEM[2585] <= 8'h80;
ROM_MEM[2586] <= 8'h2F;
ROM_MEM[2587] <= 8'h03;
ROM_MEM[2588] <= 8'hCC;
ROM_MEM[2589] <= 8'h01;
ROM_MEM[2590] <= 8'h80;
ROM_MEM[2591] <= 8'hE3;
ROM_MEM[2592] <= 8'h44;
ROM_MEM[2593] <= 8'hED;
ROM_MEM[2594] <= 8'h44;
ROM_MEM[2595] <= 8'h20;
ROM_MEM[2596] <= 8'h58;
ROM_MEM[2597] <= 8'hEE;
ROM_MEM[2598] <= 8'h84;
ROM_MEM[2599] <= 8'hCC;
ROM_MEM[2600] <= 8'hFF;
ROM_MEM[2601] <= 8'h00;
ROM_MEM[2602] <= 8'hE3;
ROM_MEM[2603] <= 8'hC4;
ROM_MEM[2604] <= 8'hED;
ROM_MEM[2605] <= 8'hC4;
ROM_MEM[2606] <= 8'hCC;
ROM_MEM[2607] <= 8'hFF;
ROM_MEM[2608] <= 8'h00;
ROM_MEM[2609] <= 8'hE3;
ROM_MEM[2610] <= 8'h42;
ROM_MEM[2611] <= 8'hED;
ROM_MEM[2612] <= 8'h42;
ROM_MEM[2613] <= 8'hFC;
ROM_MEM[2614] <= 8'h50;
ROM_MEM[2615] <= 8'h9C;
ROM_MEM[2616] <= 8'hC3;
ROM_MEM[2617] <= 8'h00;
ROM_MEM[2618] <= 8'h80;
ROM_MEM[2619] <= 8'hA3;
ROM_MEM[2620] <= 8'h44;
ROM_MEM[2621] <= 8'h2B;
ROM_MEM[2622] <= 8'h10;
ROM_MEM[2623] <= 8'hBD;
ROM_MEM[2624] <= 8'hCD;
ROM_MEM[2625] <= 8'hA2;
ROM_MEM[2626] <= 8'h10;
ROM_MEM[2627] <= 8'h83;
ROM_MEM[2628] <= 8'h01;
ROM_MEM[2629] <= 8'h80;
ROM_MEM[2630] <= 8'h2F;
ROM_MEM[2631] <= 8'h03;
ROM_MEM[2632] <= 8'hCC;
ROM_MEM[2633] <= 8'h01;
ROM_MEM[2634] <= 8'h80;
ROM_MEM[2635] <= 8'hE3;
ROM_MEM[2636] <= 8'h44;
ROM_MEM[2637] <= 8'hED;
ROM_MEM[2638] <= 8'h44;
ROM_MEM[2639] <= 8'h20;
ROM_MEM[2640] <= 8'h2C;
ROM_MEM[2641] <= 8'hEE;
ROM_MEM[2642] <= 8'h84;
ROM_MEM[2643] <= 8'hCC;
ROM_MEM[2644] <= 8'hFF;
ROM_MEM[2645] <= 8'h00;
ROM_MEM[2646] <= 8'hE3;
ROM_MEM[2647] <= 8'hC4;
ROM_MEM[2648] <= 8'hED;
ROM_MEM[2649] <= 8'hC4;
ROM_MEM[2650] <= 8'hCC;
ROM_MEM[2651] <= 8'h01;
ROM_MEM[2652] <= 8'h00;
ROM_MEM[2653] <= 8'hE3;
ROM_MEM[2654] <= 8'h42;
ROM_MEM[2655] <= 8'hED;
ROM_MEM[2656] <= 8'h42;
ROM_MEM[2657] <= 8'hFC;
ROM_MEM[2658] <= 8'h50;
ROM_MEM[2659] <= 8'h9C;
ROM_MEM[2660] <= 8'hC3;
ROM_MEM[2661] <= 8'h00;
ROM_MEM[2662] <= 8'h80;
ROM_MEM[2663] <= 8'hA3;
ROM_MEM[2664] <= 8'h44;
ROM_MEM[2665] <= 8'h2B;
ROM_MEM[2666] <= 8'h10;
ROM_MEM[2667] <= 8'hBD;
ROM_MEM[2668] <= 8'hCD;
ROM_MEM[2669] <= 8'hA2;
ROM_MEM[2670] <= 8'h10;
ROM_MEM[2671] <= 8'h83;
ROM_MEM[2672] <= 8'h01;
ROM_MEM[2673] <= 8'h80;
ROM_MEM[2674] <= 8'h2F;
ROM_MEM[2675] <= 8'h03;
ROM_MEM[2676] <= 8'hCC;
ROM_MEM[2677] <= 8'h01;
ROM_MEM[2678] <= 8'h80;
ROM_MEM[2679] <= 8'hE3;
ROM_MEM[2680] <= 8'h44;
ROM_MEM[2681] <= 8'hED;
ROM_MEM[2682] <= 8'h44;
ROM_MEM[2683] <= 8'h20;
ROM_MEM[2684] <= 8'h00;
ROM_MEM[2685] <= 8'hA6;
ROM_MEM[2686] <= 8'h03;
ROM_MEM[2687] <= 8'h85;
ROM_MEM[2688] <= 8'h02;
ROM_MEM[2689] <= 8'h27;
ROM_MEM[2690] <= 8'h02;
ROM_MEM[2691] <= 8'h6F;
ROM_MEM[2692] <= 8'h03;
ROM_MEM[2693] <= 8'h39;
ROM_MEM[2694] <= 8'hEE;
ROM_MEM[2695] <= 8'h84;
ROM_MEM[2696] <= 8'hBD;
ROM_MEM[2697] <= 8'hA9;
ROM_MEM[2698] <= 8'h0C;
ROM_MEM[2699] <= 8'hFC;
ROM_MEM[2700] <= 8'h50;
ROM_MEM[2701] <= 8'h9C;
ROM_MEM[2702] <= 8'hA3;
ROM_MEM[2703] <= 8'h44;
ROM_MEM[2704] <= 8'h2B;
ROM_MEM[2705] <= 8'h07;
ROM_MEM[2706] <= 8'hBD;
ROM_MEM[2707] <= 8'hCD;
ROM_MEM[2708] <= 8'hA0;
ROM_MEM[2709] <= 8'hE3;
ROM_MEM[2710] <= 8'h44;
ROM_MEM[2711] <= 8'hED;
ROM_MEM[2712] <= 8'h44;
ROM_MEM[2713] <= 8'hB6;
ROM_MEM[2714] <= 8'h4B;
ROM_MEM[2715] <= 8'h19;
ROM_MEM[2716] <= 8'h81;
ROM_MEM[2717] <= 8'h01;
ROM_MEM[2718] <= 8'h25;
ROM_MEM[2719] <= 8'h05;
ROM_MEM[2720] <= 8'hFC;
ROM_MEM[2721] <= 8'h50;
ROM_MEM[2722] <= 8'h9A;
ROM_MEM[2723] <= 8'h20;
ROM_MEM[2724] <= 8'h03;
ROM_MEM[2725] <= 8'hCC;
ROM_MEM[2726] <= 8'hFE;
ROM_MEM[2727] <= 8'h80;
ROM_MEM[2728] <= 8'hA3;
ROM_MEM[2729] <= 8'h42;
ROM_MEM[2730] <= 8'h2B;
ROM_MEM[2731] <= 8'h07;
ROM_MEM[2732] <= 8'hBD;
ROM_MEM[2733] <= 8'hCD;
ROM_MEM[2734] <= 8'hA0;
ROM_MEM[2735] <= 8'hE3;
ROM_MEM[2736] <= 8'h42;
ROM_MEM[2737] <= 8'hED;
ROM_MEM[2738] <= 8'h42;
ROM_MEM[2739] <= 8'h20;
ROM_MEM[2740] <= 8'hC8;
ROM_MEM[2741] <= 8'hEE;
ROM_MEM[2742] <= 8'h84;
ROM_MEM[2743] <= 8'hBD;
ROM_MEM[2744] <= 8'hA9;
ROM_MEM[2745] <= 8'h0C;
ROM_MEM[2746] <= 8'hFC;
ROM_MEM[2747] <= 8'h50;
ROM_MEM[2748] <= 8'h9C;
ROM_MEM[2749] <= 8'hA3;
ROM_MEM[2750] <= 8'h44;
ROM_MEM[2751] <= 8'h2B;
ROM_MEM[2752] <= 8'h07;
ROM_MEM[2753] <= 8'hBD;
ROM_MEM[2754] <= 8'hCD;
ROM_MEM[2755] <= 8'hA0;
ROM_MEM[2756] <= 8'hE3;
ROM_MEM[2757] <= 8'h44;
ROM_MEM[2758] <= 8'hED;
ROM_MEM[2759] <= 8'h44;
ROM_MEM[2760] <= 8'hB6;
ROM_MEM[2761] <= 8'h4B;
ROM_MEM[2762] <= 8'h19;
ROM_MEM[2763] <= 8'h81;
ROM_MEM[2764] <= 8'h01;
ROM_MEM[2765] <= 8'h25;
ROM_MEM[2766] <= 8'h05;
ROM_MEM[2767] <= 8'hFC;
ROM_MEM[2768] <= 8'h50;
ROM_MEM[2769] <= 8'h9A;
ROM_MEM[2770] <= 8'h20;
ROM_MEM[2771] <= 8'h03;
ROM_MEM[2772] <= 8'hCC;
ROM_MEM[2773] <= 8'h01;
ROM_MEM[2774] <= 8'h80;
ROM_MEM[2775] <= 8'hA3;
ROM_MEM[2776] <= 8'h42;
ROM_MEM[2777] <= 8'h2A;
ROM_MEM[2778] <= 8'h07;
ROM_MEM[2779] <= 8'hBD;
ROM_MEM[2780] <= 8'hCD;
ROM_MEM[2781] <= 8'hA0;
ROM_MEM[2782] <= 8'hE3;
ROM_MEM[2783] <= 8'h42;
ROM_MEM[2784] <= 8'hED;
ROM_MEM[2785] <= 8'h42;
ROM_MEM[2786] <= 8'h20;
ROM_MEM[2787] <= 8'h99;
ROM_MEM[2788] <= 8'h8E;
ROM_MEM[2789] <= 8'h49;
ROM_MEM[2790] <= 8'h4B;
ROM_MEM[2791] <= 8'h9F;
ROM_MEM[2792] <= 8'hA8;
ROM_MEM[2793] <= 8'hA6;
ROM_MEM[2794] <= 8'h03;
ROM_MEM[2795] <= 8'h10;
ROM_MEM[2796] <= 8'h27;
ROM_MEM[2797] <= 8'h01;
ROM_MEM[2798] <= 8'h45;
ROM_MEM[2799] <= 8'h85;
ROM_MEM[2800] <= 8'h10;
ROM_MEM[2801] <= 8'h27;
ROM_MEM[2802] <= 8'h06;
ROM_MEM[2803] <= 8'hBD;
ROM_MEM[2804] <= 8'hAC;
ROM_MEM[2805] <= 8'hB1;
ROM_MEM[2806] <= 8'h7E;
ROM_MEM[2807] <= 8'hAC;
ROM_MEM[2808] <= 8'h34;
ROM_MEM[2809] <= 8'h85;
ROM_MEM[2810] <= 8'h04;
ROM_MEM[2811] <= 8'h27;
ROM_MEM[2812] <= 8'h14;
ROM_MEM[2813] <= 8'hFC;
ROM_MEM[2814] <= 8'h50;
ROM_MEM[2815] <= 8'h98;
ROM_MEM[2816] <= 8'hFD;
ROM_MEM[2817] <= 8'h50;
ROM_MEM[2818] <= 8'h40;
ROM_MEM[2819] <= 8'hFC;
ROM_MEM[2820] <= 8'h50;
ROM_MEM[2821] <= 8'h9A;
ROM_MEM[2822] <= 8'hFD;
ROM_MEM[2823] <= 8'h50;
ROM_MEM[2824] <= 8'h42;
ROM_MEM[2825] <= 8'hFC;
ROM_MEM[2826] <= 8'h50;
ROM_MEM[2827] <= 8'h9C;
ROM_MEM[2828] <= 8'hFD;
ROM_MEM[2829] <= 8'h50;
ROM_MEM[2830] <= 8'h44;
ROM_MEM[2831] <= 8'h20;
ROM_MEM[2832] <= 8'h0C;
ROM_MEM[2833] <= 8'hCC;
ROM_MEM[2834] <= 8'h00;
ROM_MEM[2835] <= 8'h00;
ROM_MEM[2836] <= 8'hFD;
ROM_MEM[2837] <= 8'h50;
ROM_MEM[2838] <= 8'h40;
ROM_MEM[2839] <= 8'hFD;
ROM_MEM[2840] <= 8'h50;
ROM_MEM[2841] <= 8'h42;
ROM_MEM[2842] <= 8'hFD;
ROM_MEM[2843] <= 8'h50;
ROM_MEM[2844] <= 8'h44;
ROM_MEM[2845] <= 8'h4F;
ROM_MEM[2846] <= 8'hE6;
ROM_MEM[2847] <= 8'h02;
ROM_MEM[2848] <= 8'hFD;
ROM_MEM[2849] <= 8'h47;
ROM_MEM[2850] <= 8'h01;
ROM_MEM[2851] <= 8'h86;
ROM_MEM[2852] <= 8'h67;
ROM_MEM[2853] <= 8'hBD;
ROM_MEM[2854] <= 8'hCD;
ROM_MEM[2855] <= 8'hBA;
ROM_MEM[2856] <= 8'hFC;
ROM_MEM[2857] <= 8'h50;
ROM_MEM[2858] <= 8'h00;
ROM_MEM[2859] <= 8'h10;
ROM_MEM[2860] <= 8'h83;
ROM_MEM[2861] <= 8'h00;
ROM_MEM[2862] <= 8'h01;
ROM_MEM[2863] <= 8'h10;
ROM_MEM[2864] <= 8'h2F;
ROM_MEM[2865] <= 8'h00;
ROM_MEM[2866] <= 8'hF4;
ROM_MEM[2867] <= 8'h10;
ROM_MEM[2868] <= 8'h83;
ROM_MEM[2869] <= 8'h7F;
ROM_MEM[2870] <= 8'h00;
ROM_MEM[2871] <= 8'h10;
ROM_MEM[2872] <= 8'h22;
ROM_MEM[2873] <= 8'h00;
ROM_MEM[2874] <= 8'hEC;
ROM_MEM[2875] <= 8'hFD;
ROM_MEM[2876] <= 8'h47;
ROM_MEM[2877] <= 8'h04;
ROM_MEM[2878] <= 8'hFD;
ROM_MEM[2879] <= 8'h50;
ROM_MEM[2880] <= 8'h18;
ROM_MEM[2881] <= 8'hFC;
ROM_MEM[2882] <= 8'h50;
ROM_MEM[2883] <= 8'h02;
ROM_MEM[2884] <= 8'hFD;
ROM_MEM[2885] <= 8'h50;
ROM_MEM[2886] <= 8'h1A;
ROM_MEM[2887] <= 8'h2A;
ROM_MEM[2888] <= 8'h04;
ROM_MEM[2889] <= 8'h43;
ROM_MEM[2890] <= 8'h50;
ROM_MEM[2891] <= 8'h82;
ROM_MEM[2892] <= 8'hFF;
ROM_MEM[2893] <= 8'hB3;
ROM_MEM[2894] <= 8'h50;
ROM_MEM[2895] <= 8'h00;
ROM_MEM[2896] <= 8'h10;
ROM_MEM[2897] <= 8'h24;
ROM_MEM[2898] <= 8'h00;
ROM_MEM[2899] <= 8'hD3;
ROM_MEM[2900] <= 8'hFC;
ROM_MEM[2901] <= 8'h50;
ROM_MEM[2902] <= 8'h04;
ROM_MEM[2903] <= 8'hFD;
ROM_MEM[2904] <= 8'h50;
ROM_MEM[2905] <= 8'h1C;
ROM_MEM[2906] <= 8'h2A;
ROM_MEM[2907] <= 8'h04;
ROM_MEM[2908] <= 8'h43;
ROM_MEM[2909] <= 8'h50;
ROM_MEM[2910] <= 8'h82;
ROM_MEM[2911] <= 8'hFF;
ROM_MEM[2912] <= 8'hB3;
ROM_MEM[2913] <= 8'h50;
ROM_MEM[2914] <= 8'h00;
ROM_MEM[2915] <= 8'h10;
ROM_MEM[2916] <= 8'h24;
ROM_MEM[2917] <= 8'h00;
ROM_MEM[2918] <= 8'hC0;
ROM_MEM[2919] <= 8'hBD;
ROM_MEM[2920] <= 8'hCC;
ROM_MEM[2921] <= 8'hF0;
ROM_MEM[2922] <= 8'h9E;
ROM_MEM[2923] <= 8'hA8;
ROM_MEM[2924] <= 8'hA6;
ROM_MEM[2925] <= 8'h03;
ROM_MEM[2926] <= 8'h85;
ROM_MEM[2927] <= 8'h03;
ROM_MEM[2928] <= 8'h27;
ROM_MEM[2929] <= 8'h4E;
ROM_MEM[2930] <= 8'hCC;
ROM_MEM[2931] <= 8'h00;
ROM_MEM[2932] <= 8'h80;
ROM_MEM[2933] <= 8'hFD;
ROM_MEM[2934] <= 8'h50;
ROM_MEM[2935] <= 8'h02;
ROM_MEM[2936] <= 8'h86;
ROM_MEM[2937] <= 8'h86;
ROM_MEM[2938] <= 8'hBD;
ROM_MEM[2939] <= 8'hCD;
ROM_MEM[2940] <= 8'hBA;
ROM_MEM[2941] <= 8'hFC;
ROM_MEM[2942] <= 8'h50;
ROM_MEM[2943] <= 8'h02;
ROM_MEM[2944] <= 8'hC3;
ROM_MEM[2945] <= 8'h00;
ROM_MEM[2946] <= 8'h0A;
ROM_MEM[2947] <= 8'hDD;
ROM_MEM[2948] <= 8'h03;
ROM_MEM[2949] <= 8'hDC;
ROM_MEM[2950] <= 8'hD6;
ROM_MEM[2951] <= 8'h93;
ROM_MEM[2952] <= 8'hB3;
ROM_MEM[2953] <= 8'h2A;
ROM_MEM[2954] <= 8'h04;
ROM_MEM[2955] <= 8'h43;
ROM_MEM[2956] <= 8'h50;
ROM_MEM[2957] <= 8'h82;
ROM_MEM[2958] <= 8'hFF;
ROM_MEM[2959] <= 8'hDD;
ROM_MEM[2960] <= 8'h01;
ROM_MEM[2961] <= 8'h93;
ROM_MEM[2962] <= 8'h03;
ROM_MEM[2963] <= 8'h2E;
ROM_MEM[2964] <= 8'h2B;
ROM_MEM[2965] <= 8'hDC;
ROM_MEM[2966] <= 8'hD8;
ROM_MEM[2967] <= 8'h93;
ROM_MEM[2968] <= 8'hB5;
ROM_MEM[2969] <= 8'h2A;
ROM_MEM[2970] <= 8'h04;
ROM_MEM[2971] <= 8'h43;
ROM_MEM[2972] <= 8'h50;
ROM_MEM[2973] <= 8'h82;
ROM_MEM[2974] <= 8'hFF;
ROM_MEM[2975] <= 8'h10;
ROM_MEM[2976] <= 8'h93;
ROM_MEM[2977] <= 8'h03;
ROM_MEM[2978] <= 8'h2E;
ROM_MEM[2979] <= 8'h1C;
ROM_MEM[2980] <= 8'hD3;
ROM_MEM[2981] <= 8'h01;
ROM_MEM[2982] <= 8'hDD;
ROM_MEM[2983] <= 8'h01;
ROM_MEM[2984] <= 8'hDC;
ROM_MEM[2985] <= 8'h03;
ROM_MEM[2986] <= 8'h44;
ROM_MEM[2987] <= 8'h56;
ROM_MEM[2988] <= 8'hD3;
ROM_MEM[2989] <= 8'h03;
ROM_MEM[2990] <= 8'h93;
ROM_MEM[2991] <= 8'h01;
ROM_MEM[2992] <= 8'h2D;
ROM_MEM[2993] <= 8'h0E;
ROM_MEM[2994] <= 8'hFC;
ROM_MEM[2995] <= 8'h50;
ROM_MEM[2996] <= 8'h18;
ROM_MEM[2997] <= 8'h10;
ROM_MEM[2998] <= 8'h93;
ROM_MEM[2999] <= 8'hCC;
ROM_MEM[3000] <= 8'h24;
ROM_MEM[3001] <= 8'h06;
ROM_MEM[3002] <= 8'hDD;
ROM_MEM[3003] <= 8'hCC;
ROM_MEM[3004] <= 8'h9E;
ROM_MEM[3005] <= 8'hA8;
ROM_MEM[3006] <= 8'h9F;
ROM_MEM[3007] <= 8'hCA;
ROM_MEM[3008] <= 8'hA6;
ROM_MEM[3009] <= 8'h03;
ROM_MEM[3010] <= 8'h85;
ROM_MEM[3011] <= 8'h01;
ROM_MEM[3012] <= 8'h27;
ROM_MEM[3013] <= 8'h5C;
ROM_MEM[3014] <= 8'hFC;
ROM_MEM[3015] <= 8'h50;
ROM_MEM[3016] <= 8'h18;
ROM_MEM[3017] <= 8'h58;
ROM_MEM[3018] <= 8'h49;
ROM_MEM[3019] <= 8'h2B;
ROM_MEM[3020] <= 8'h55;
ROM_MEM[3021] <= 8'hFE;
ROM_MEM[3022] <= 8'h50;
ROM_MEM[3023] <= 8'h86;
ROM_MEM[3024] <= 8'h11;
ROM_MEM[3025] <= 8'h83;
ROM_MEM[3026] <= 8'h02;
ROM_MEM[3027] <= 8'h00;
ROM_MEM[3028] <= 8'h2D;
ROM_MEM[3029] <= 8'h05;
ROM_MEM[3030] <= 8'hB3;
ROM_MEM[3031] <= 8'h50;
ROM_MEM[3032] <= 8'h86;
ROM_MEM[3033] <= 8'h20;
ROM_MEM[3034] <= 8'h03;
ROM_MEM[3035] <= 8'h83;
ROM_MEM[3036] <= 8'h02;
ROM_MEM[3037] <= 8'h00;
ROM_MEM[3038] <= 8'h2F;
ROM_MEM[3039] <= 8'h05;
ROM_MEM[3040] <= 8'h83;
ROM_MEM[3041] <= 8'h01;
ROM_MEM[3042] <= 8'h10;
ROM_MEM[3043] <= 8'h2E;
ROM_MEM[3044] <= 8'h3D;
ROM_MEM[3045] <= 8'hDC;
ROM_MEM[3046] <= 8'hD6;
ROM_MEM[3047] <= 8'h2B;
ROM_MEM[3048] <= 8'h07;
ROM_MEM[3049] <= 8'h83;
ROM_MEM[3050] <= 8'h01;
ROM_MEM[3051] <= 8'hC0;
ROM_MEM[3052] <= 8'h2C;
ROM_MEM[3053] <= 8'h34;
ROM_MEM[3054] <= 8'h20;
ROM_MEM[3055] <= 8'h05;
ROM_MEM[3056] <= 8'h83;
ROM_MEM[3057] <= 8'hFE;
ROM_MEM[3058] <= 8'h40;
ROM_MEM[3059] <= 8'h2F;
ROM_MEM[3060] <= 8'h2D;
ROM_MEM[3061] <= 8'hDC;
ROM_MEM[3062] <= 8'hD8;
ROM_MEM[3063] <= 8'h2B;
ROM_MEM[3064] <= 8'h07;
ROM_MEM[3065] <= 8'h83;
ROM_MEM[3066] <= 8'h01;
ROM_MEM[3067] <= 8'hE0;
ROM_MEM[3068] <= 8'h2C;
ROM_MEM[3069] <= 8'h24;
ROM_MEM[3070] <= 8'h20;
ROM_MEM[3071] <= 8'h05;
ROM_MEM[3072] <= 8'h83;
ROM_MEM[3073] <= 8'hFE;
ROM_MEM[3074] <= 8'h60;
ROM_MEM[3075] <= 8'h2F;
ROM_MEM[3076] <= 8'h1D;
ROM_MEM[3077] <= 8'h9C;
ROM_MEM[3078] <= 8'hCA;
ROM_MEM[3079] <= 8'h26;
ROM_MEM[3080] <= 8'h0B;
ROM_MEM[3081] <= 8'h96;
ROM_MEM[3082] <= 8'hBC;
ROM_MEM[3083] <= 8'h27;
ROM_MEM[3084] <= 8'h07;
ROM_MEM[3085] <= 8'hBD;
ROM_MEM[3086] <= 8'hAD;
ROM_MEM[3087] <= 8'h20;
ROM_MEM[3088] <= 8'h9E;
ROM_MEM[3089] <= 8'hA8;
ROM_MEM[3090] <= 8'h20;
ROM_MEM[3091] <= 8'h0E;
ROM_MEM[3092] <= 8'hBD;
ROM_MEM[3093] <= 8'hAC;
ROM_MEM[3094] <= 8'hE0;
ROM_MEM[3095] <= 8'hCC;
ROM_MEM[3096] <= 8'h80;
ROM_MEM[3097] <= 8'h40;
ROM_MEM[3098] <= 8'hED;
ROM_MEM[3099] <= 8'hA1;
ROM_MEM[3100] <= 8'hBD;
ROM_MEM[3101] <= 8'hAC;
ROM_MEM[3102] <= 8'hB1;
ROM_MEM[3103] <= 8'h7E;
ROM_MEM[3104] <= 8'hAC;
ROM_MEM[3105] <= 8'h34;
ROM_MEM[3106] <= 8'hBD;
ROM_MEM[3107] <= 8'hAC;
ROM_MEM[3108] <= 8'h52;
ROM_MEM[3109] <= 8'h20;
ROM_MEM[3110] <= 8'h0D;
ROM_MEM[3111] <= 8'hA6;
ROM_MEM[3112] <= 8'h03;
ROM_MEM[3113] <= 8'h85;
ROM_MEM[3114] <= 8'h01;
ROM_MEM[3115] <= 8'h27;
ROM_MEM[3116] <= 8'h04;
ROM_MEM[3117] <= 8'h86;
ROM_MEM[3118] <= 8'h00;
ROM_MEM[3119] <= 8'h20;
ROM_MEM[3120] <= 8'h01;
ROM_MEM[3121] <= 8'h4F;
ROM_MEM[3122] <= 8'hA7;
ROM_MEM[3123] <= 8'h03;
ROM_MEM[3124] <= 8'h9E;
ROM_MEM[3125] <= 8'hA8;
ROM_MEM[3126] <= 8'h30;
ROM_MEM[3127] <= 8'h06;
ROM_MEM[3128] <= 8'h8C;
ROM_MEM[3129] <= 8'h49;
ROM_MEM[3130] <= 8'h6F;
ROM_MEM[3131] <= 8'h10;
ROM_MEM[3132] <= 8'h25;
ROM_MEM[3133] <= 8'hFE;
ROM_MEM[3134] <= 8'hA8;
ROM_MEM[3135] <= 8'hFC;
ROM_MEM[3136] <= 8'h50;
ROM_MEM[3137] <= 8'h98;
ROM_MEM[3138] <= 8'hFD;
ROM_MEM[3139] <= 8'h50;
ROM_MEM[3140] <= 8'h40;
ROM_MEM[3141] <= 8'hFC;
ROM_MEM[3142] <= 8'h50;
ROM_MEM[3143] <= 8'h9A;
ROM_MEM[3144] <= 8'hFD;
ROM_MEM[3145] <= 8'h50;
ROM_MEM[3146] <= 8'h42;
ROM_MEM[3147] <= 8'hFC;
ROM_MEM[3148] <= 8'h50;
ROM_MEM[3149] <= 8'h9C;
ROM_MEM[3150] <= 8'hFD;
ROM_MEM[3151] <= 8'h50;
ROM_MEM[3152] <= 8'h44;
ROM_MEM[3153] <= 8'h39;
ROM_MEM[3154] <= 8'h9E;
ROM_MEM[3155] <= 8'hA8;
ROM_MEM[3156] <= 8'h86;
ROM_MEM[3157] <= 8'h08;
ROM_MEM[3158] <= 8'h97;
ROM_MEM[3159] <= 8'h01;
ROM_MEM[3160] <= 8'hFC;
ROM_MEM[3161] <= 8'h50;
ROM_MEM[3162] <= 8'h18;
ROM_MEM[3163] <= 8'h0A;
ROM_MEM[3164] <= 8'h01;
ROM_MEM[3165] <= 8'h27;
ROM_MEM[3166] <= 8'h06;
ROM_MEM[3167] <= 8'h58;
ROM_MEM[3168] <= 8'h49;
ROM_MEM[3169] <= 8'h2A;
ROM_MEM[3170] <= 8'hF8;
ROM_MEM[3171] <= 8'h84;
ROM_MEM[3172] <= 8'h7F;
ROM_MEM[3173] <= 8'h97;
ROM_MEM[3174] <= 8'h02;
ROM_MEM[3175] <= 8'hA6;
ROM_MEM[3176] <= 8'h03;
ROM_MEM[3177] <= 8'h84;
ROM_MEM[3178] <= 8'h20;
ROM_MEM[3179] <= 8'h26;
ROM_MEM[3180] <= 8'h0F;
ROM_MEM[3181] <= 8'h96;
ROM_MEM[3182] <= 8'h01;
ROM_MEM[3183] <= 8'h8A;
ROM_MEM[3184] <= 8'h70;
ROM_MEM[3185] <= 8'hD6;
ROM_MEM[3186] <= 8'h02;
ROM_MEM[3187] <= 8'hED;
ROM_MEM[3188] <= 8'hA1;
ROM_MEM[3189] <= 8'hCC;
ROM_MEM[3190] <= 8'hA0;
ROM_MEM[3191] <= 8'h15;
ROM_MEM[3192] <= 8'hED;
ROM_MEM[3193] <= 8'hA1;
ROM_MEM[3194] <= 8'h20;
ROM_MEM[3195] <= 8'h2A;
ROM_MEM[3196] <= 8'hD6;
ROM_MEM[3197] <= 8'h02;
ROM_MEM[3198] <= 8'h96;
ROM_MEM[3199] <= 8'h01;
ROM_MEM[3200] <= 8'h4C;
ROM_MEM[3201] <= 8'h81;
ROM_MEM[3202] <= 8'h03;
ROM_MEM[3203] <= 8'h24;
ROM_MEM[3204] <= 8'h05;
ROM_MEM[3205] <= 8'h86;
ROM_MEM[3206] <= 8'h03;
ROM_MEM[3207] <= 8'h5F;
ROM_MEM[3208] <= 8'h20;
ROM_MEM[3209] <= 8'h07;
ROM_MEM[3210] <= 8'h81;
ROM_MEM[3211] <= 8'h06;
ROM_MEM[3212] <= 8'h25;
ROM_MEM[3213] <= 8'h03;
ROM_MEM[3214] <= 8'h86;
ROM_MEM[3215] <= 8'h06;
ROM_MEM[3216] <= 8'h5F;
ROM_MEM[3217] <= 8'h8A;
ROM_MEM[3218] <= 8'h70;
ROM_MEM[3219] <= 8'hED;
ROM_MEM[3220] <= 8'hA1;
ROM_MEM[3221] <= 8'hE6;
ROM_MEM[3222] <= 8'h05;
ROM_MEM[3223] <= 8'h58;
ROM_MEM[3224] <= 8'h58;
ROM_MEM[3225] <= 8'h58;
ROM_MEM[3226] <= 8'h58;
ROM_MEM[3227] <= 8'hCA;
ROM_MEM[3228] <= 8'h0F;
ROM_MEM[3229] <= 8'h86;
ROM_MEM[3230] <= 8'h65;
ROM_MEM[3231] <= 8'hED;
ROM_MEM[3232] <= 8'hA1;
ROM_MEM[3233] <= 8'hCC;
ROM_MEM[3234] <= 8'hA0;
ROM_MEM[3235] <= 8'h17;
ROM_MEM[3236] <= 8'hED;
ROM_MEM[3237] <= 8'hA1;
ROM_MEM[3238] <= 8'hCC;
ROM_MEM[3239] <= 8'h72;
ROM_MEM[3240] <= 8'h00;
ROM_MEM[3241] <= 8'hED;
ROM_MEM[3242] <= 8'hA1;
ROM_MEM[3243] <= 8'hCC;
ROM_MEM[3244] <= 8'h80;
ROM_MEM[3245] <= 8'h40;
ROM_MEM[3246] <= 8'hED;
ROM_MEM[3247] <= 8'hA1;
ROM_MEM[3248] <= 8'h39;
ROM_MEM[3249] <= 8'h9E;
ROM_MEM[3250] <= 8'hA8;
ROM_MEM[3251] <= 8'hEE;
ROM_MEM[3252] <= 8'h84;
ROM_MEM[3253] <= 8'hEC;
ROM_MEM[3254] <= 8'hC4;
ROM_MEM[3255] <= 8'hED;
ROM_MEM[3256] <= 8'hA1;
ROM_MEM[3257] <= 8'hEC;
ROM_MEM[3258] <= 8'h42;
ROM_MEM[3259] <= 8'hED;
ROM_MEM[3260] <= 8'hA1;
ROM_MEM[3261] <= 8'hA6;
ROM_MEM[3262] <= 8'h05;
ROM_MEM[3263] <= 8'hC6;
ROM_MEM[3264] <= 8'h10;
ROM_MEM[3265] <= 8'h3D;
ROM_MEM[3266] <= 8'h86;
ROM_MEM[3267] <= 8'h70;
ROM_MEM[3268] <= 8'hED;
ROM_MEM[3269] <= 8'hA1;
ROM_MEM[3270] <= 8'hE6;
ROM_MEM[3271] <= 8'h05;
ROM_MEM[3272] <= 8'h58;
ROM_MEM[3273] <= 8'h58;
ROM_MEM[3274] <= 8'h58;
ROM_MEM[3275] <= 8'h58;
ROM_MEM[3276] <= 8'h86;
ROM_MEM[3277] <= 8'h67;
ROM_MEM[3278] <= 8'hED;
ROM_MEM[3279] <= 8'hA1;
ROM_MEM[3280] <= 8'hCC;
ROM_MEM[3281] <= 8'hA0;
ROM_MEM[3282] <= 8'h17;
ROM_MEM[3283] <= 8'hED;
ROM_MEM[3284] <= 8'hA1;
ROM_MEM[3285] <= 8'hCC;
ROM_MEM[3286] <= 8'h72;
ROM_MEM[3287] <= 8'h00;
ROM_MEM[3288] <= 8'hED;
ROM_MEM[3289] <= 8'hA1;
ROM_MEM[3290] <= 8'hCC;
ROM_MEM[3291] <= 8'h80;
ROM_MEM[3292] <= 8'h40;
ROM_MEM[3293] <= 8'hED;
ROM_MEM[3294] <= 8'hA1;
ROM_MEM[3295] <= 8'h39;
ROM_MEM[3296] <= 8'hEE;
ROM_MEM[3297] <= 8'h84;
ROM_MEM[3298] <= 8'hEC;
ROM_MEM[3299] <= 8'h3C;
ROM_MEM[3300] <= 8'hED;
ROM_MEM[3301] <= 8'hC4;
ROM_MEM[3302] <= 8'hEC;
ROM_MEM[3303] <= 8'h3E;
ROM_MEM[3304] <= 8'hED;
ROM_MEM[3305] <= 8'h42;
ROM_MEM[3306] <= 8'h86;
ROM_MEM[3307] <= 8'h10;
ROM_MEM[3308] <= 8'hA7;
ROM_MEM[3309] <= 8'h03;
ROM_MEM[3310] <= 8'h86;
ROM_MEM[3311] <= 8'h0F;
ROM_MEM[3312] <= 8'hA7;
ROM_MEM[3313] <= 8'h05;
ROM_MEM[3314] <= 8'h86;
ROM_MEM[3315] <= 8'h00;
ROM_MEM[3316] <= 8'hA7;
ROM_MEM[3317] <= 8'h04;
ROM_MEM[3318] <= 8'hBD;
ROM_MEM[3319] <= 8'h98;
ROM_MEM[3320] <= 8'h74;
ROM_MEM[3321] <= 8'h96;
ROM_MEM[3322] <= 8'h63;
ROM_MEM[3323] <= 8'h26;
ROM_MEM[3324] <= 8'h03;
ROM_MEM[3325] <= 8'hB6;
ROM_MEM[3326] <= 8'h47;
ROM_MEM[3327] <= 8'h03;
ROM_MEM[3328] <= 8'hC6;
ROM_MEM[3329] <= 8'h20;
ROM_MEM[3330] <= 8'h4D;
ROM_MEM[3331] <= 8'h2A;
ROM_MEM[3332] <= 8'h01;
ROM_MEM[3333] <= 8'h50;
ROM_MEM[3334] <= 8'hD7;
ROM_MEM[3335] <= 8'h63;
ROM_MEM[3336] <= 8'hBD;
ROM_MEM[3337] <= 8'hBD;
ROM_MEM[3338] <= 8'hF3;
ROM_MEM[3339] <= 8'hB6;
ROM_MEM[3340] <= 8'h4B;
ROM_MEM[3341] <= 8'h37;
ROM_MEM[3342] <= 8'h26;
ROM_MEM[3343] <= 8'h0F;
ROM_MEM[3344] <= 8'h7C;
ROM_MEM[3345] <= 8'h4B;
ROM_MEM[3346] <= 8'h37;
ROM_MEM[3347] <= 8'h96;
ROM_MEM[3348] <= 8'h60;
ROM_MEM[3349] <= 8'h81;
ROM_MEM[3350] <= 8'h03;
ROM_MEM[3351] <= 8'h23;
ROM_MEM[3352] <= 8'h06;
ROM_MEM[3353] <= 8'hBD;
ROM_MEM[3354] <= 8'hBD;
ROM_MEM[3355] <= 8'h21;
ROM_MEM[3356] <= 8'hBD;
ROM_MEM[3357] <= 8'hBD;
ROM_MEM[3358] <= 8'hE9;
ROM_MEM[3359] <= 8'h39;
ROM_MEM[3360] <= 8'hDE;
ROM_MEM[3361] <= 8'hCA;
ROM_MEM[3362] <= 8'hA6;
ROM_MEM[3363] <= 8'h43;
ROM_MEM[3364] <= 8'h27;
ROM_MEM[3365] <= 8'h17;
ROM_MEM[3366] <= 8'h84;
ROM_MEM[3367] <= 8'h04;
ROM_MEM[3368] <= 8'h8A;
ROM_MEM[3369] <= 8'h20;
ROM_MEM[3370] <= 8'hA7;
ROM_MEM[3371] <= 8'h43;
ROM_MEM[3372] <= 8'h86;
ROM_MEM[3373] <= 8'h0F;
ROM_MEM[3374] <= 8'hA7;
ROM_MEM[3375] <= 8'h45;
ROM_MEM[3376] <= 8'h86;
ROM_MEM[3377] <= 8'h00;
ROM_MEM[3378] <= 8'hA7;
ROM_MEM[3379] <= 8'h44;
ROM_MEM[3380] <= 8'hBD;
ROM_MEM[3381] <= 8'hBE;
ROM_MEM[3382] <= 8'h07;
ROM_MEM[3383] <= 8'hBD;
ROM_MEM[3384] <= 8'h98;
ROM_MEM[3385] <= 8'h01;
ROM_MEM[3386] <= 8'hBD;
ROM_MEM[3387] <= 8'hBD;
ROM_MEM[3388] <= 8'hF8;
ROM_MEM[3389] <= 8'h39;
ROM_MEM[3390] <= 8'h86;
ROM_MEM[3391] <= 8'h01;
ROM_MEM[3392] <= 8'h97;
ROM_MEM[3393] <= 8'h45;
ROM_MEM[3394] <= 8'hFC;
ROM_MEM[3395] <= 8'h50;
ROM_MEM[3396] <= 8'h98;
ROM_MEM[3397] <= 8'hC3;
ROM_MEM[3398] <= 8'h01;
ROM_MEM[3399] <= 8'h00;
ROM_MEM[3400] <= 8'hDD;
ROM_MEM[3401] <= 8'h46;
ROM_MEM[3402] <= 8'hFC;
ROM_MEM[3403] <= 8'h50;
ROM_MEM[3404] <= 8'h9A;
ROM_MEM[3405] <= 8'hDD;
ROM_MEM[3406] <= 8'h48;
ROM_MEM[3407] <= 8'hFC;
ROM_MEM[3408] <= 8'h50;
ROM_MEM[3409] <= 8'h9C;
ROM_MEM[3410] <= 8'hDD;
ROM_MEM[3411] <= 8'h4A;
ROM_MEM[3412] <= 8'h8E;
ROM_MEM[3413] <= 8'h49;
ROM_MEM[3414] <= 8'h4B;
ROM_MEM[3415] <= 8'h9F;
ROM_MEM[3416] <= 8'hCA;
ROM_MEM[3417] <= 8'hBD;
ROM_MEM[3418] <= 8'hAD;
ROM_MEM[3419] <= 8'h20;
ROM_MEM[3420] <= 8'h9E;
ROM_MEM[3421] <= 8'hCA;
ROM_MEM[3422] <= 8'h30;
ROM_MEM[3423] <= 8'h06;
ROM_MEM[3424] <= 8'h8C;
ROM_MEM[3425] <= 8'h49;
ROM_MEM[3426] <= 8'h6F;
ROM_MEM[3427] <= 8'h25;
ROM_MEM[3428] <= 8'hF2;
ROM_MEM[3429] <= 8'hBD;
ROM_MEM[3430] <= 8'hBD;
ROM_MEM[3431] <= 8'hA3;
ROM_MEM[3432] <= 8'hBD;
ROM_MEM[3433] <= 8'hBD;
ROM_MEM[3434] <= 8'hD5;
ROM_MEM[3435] <= 8'h39;
ROM_MEM[3436] <= 8'h96;
ROM_MEM[3437] <= 8'h45;
ROM_MEM[3438] <= 8'h27;
ROM_MEM[3439] <= 8'h3E;
ROM_MEM[3440] <= 8'hDC;
ROM_MEM[3441] <= 8'h46;
ROM_MEM[3442] <= 8'hC3;
ROM_MEM[3443] <= 8'h03;
ROM_MEM[3444] <= 8'h00;
ROM_MEM[3445] <= 8'hF3;
ROM_MEM[3446] <= 8'h50;
ROM_MEM[3447] <= 8'h86;
ROM_MEM[3448] <= 8'h10;
ROM_MEM[3449] <= 8'h93;
ROM_MEM[3450] <= 8'h96;
ROM_MEM[3451] <= 8'h2B;
ROM_MEM[3452] <= 8'h02;
ROM_MEM[3453] <= 8'hDC;
ROM_MEM[3454] <= 8'h96;
ROM_MEM[3455] <= 8'hDD;
ROM_MEM[3456] <= 8'h46;
ROM_MEM[3457] <= 8'hDC;
ROM_MEM[3458] <= 8'h96;
ROM_MEM[3459] <= 8'h93;
ROM_MEM[3460] <= 8'h46;
ROM_MEM[3461] <= 8'h83;
ROM_MEM[3462] <= 8'h10;
ROM_MEM[3463] <= 8'h00;
ROM_MEM[3464] <= 8'h10;
ROM_MEM[3465] <= 8'h93;
ROM_MEM[3466] <= 8'h4A;
ROM_MEM[3467] <= 8'h2C;
ROM_MEM[3468] <= 8'h02;
ROM_MEM[3469] <= 8'hDD;
ROM_MEM[3470] <= 8'h4A;
ROM_MEM[3471] <= 8'hDC;
ROM_MEM[3472] <= 8'h96;
ROM_MEM[3473] <= 8'h93;
ROM_MEM[3474] <= 8'h46;
ROM_MEM[3475] <= 8'hBD;
ROM_MEM[3476] <= 8'hCD;
ROM_MEM[3477] <= 8'hA0;
ROM_MEM[3478] <= 8'h0D;
ROM_MEM[3479] <= 8'h48;
ROM_MEM[3480] <= 8'h2B;
ROM_MEM[3481] <= 8'h09;
ROM_MEM[3482] <= 8'h10;
ROM_MEM[3483] <= 8'h93;
ROM_MEM[3484] <= 8'h48;
ROM_MEM[3485] <= 8'h2C;
ROM_MEM[3486] <= 8'h02;
ROM_MEM[3487] <= 8'hDD;
ROM_MEM[3488] <= 8'h48;
ROM_MEM[3489] <= 8'h20;
ROM_MEM[3490] <= 8'h0B;
ROM_MEM[3491] <= 8'h43;
ROM_MEM[3492] <= 8'h50;
ROM_MEM[3493] <= 8'h82;
ROM_MEM[3494] <= 8'hFF;
ROM_MEM[3495] <= 8'h10;
ROM_MEM[3496] <= 8'h93;
ROM_MEM[3497] <= 8'h48;
ROM_MEM[3498] <= 8'h2F;
ROM_MEM[3499] <= 8'h02;
ROM_MEM[3500] <= 8'hDD;
ROM_MEM[3501] <= 8'h48;
ROM_MEM[3502] <= 8'h39;
ROM_MEM[3503] <= 8'h96;
ROM_MEM[3504] <= 8'h45;
ROM_MEM[3505] <= 8'h27;
ROM_MEM[3506] <= 8'h20;
ROM_MEM[3507] <= 8'hDC;
ROM_MEM[3508] <= 8'h46;
ROM_MEM[3509] <= 8'hFD;
ROM_MEM[3510] <= 8'h50;
ROM_MEM[3511] <= 8'h78;
ROM_MEM[3512] <= 8'hDC;
ROM_MEM[3513] <= 8'h48;
ROM_MEM[3514] <= 8'hC3;
ROM_MEM[3515] <= 8'h00;
ROM_MEM[3516] <= 8'h80;
ROM_MEM[3517] <= 8'hFD;
ROM_MEM[3518] <= 8'h50;
ROM_MEM[3519] <= 8'h7A;
ROM_MEM[3520] <= 8'hDC;
ROM_MEM[3521] <= 8'h4A;
ROM_MEM[3522] <= 8'hFD;
ROM_MEM[3523] <= 8'h50;
ROM_MEM[3524] <= 8'h7C;
ROM_MEM[3525] <= 8'hBD;
ROM_MEM[3526] <= 8'hAD;
ROM_MEM[3527] <= 8'hD4;
ROM_MEM[3528] <= 8'hDC;
ROM_MEM[3529] <= 8'h48;
ROM_MEM[3530] <= 8'h83;
ROM_MEM[3531] <= 8'h00;
ROM_MEM[3532] <= 8'h80;
ROM_MEM[3533] <= 8'hFD;
ROM_MEM[3534] <= 8'h50;
ROM_MEM[3535] <= 8'h7A;
ROM_MEM[3536] <= 8'hBD;
ROM_MEM[3537] <= 8'hAD;
ROM_MEM[3538] <= 8'hD4;
ROM_MEM[3539] <= 8'h39;
ROM_MEM[3540] <= 8'hCC;
ROM_MEM[3541] <= 8'h00;
ROM_MEM[3542] <= 8'h0F;
ROM_MEM[3543] <= 8'hFD;
ROM_MEM[3544] <= 8'h47;
ROM_MEM[3545] <= 8'h01;
ROM_MEM[3546] <= 8'h86;
ROM_MEM[3547] <= 8'h67;
ROM_MEM[3548] <= 8'hBD;
ROM_MEM[3549] <= 8'hCD;
ROM_MEM[3550] <= 8'hBA;
ROM_MEM[3551] <= 8'hFC;
ROM_MEM[3552] <= 8'h50;
ROM_MEM[3553] <= 8'h00;
ROM_MEM[3554] <= 8'h83;
ROM_MEM[3555] <= 8'hE0;
ROM_MEM[3556] <= 8'h00;
ROM_MEM[3557] <= 8'h2E;
ROM_MEM[3558] <= 8'h04;
ROM_MEM[3559] <= 8'h86;
ROM_MEM[3560] <= 8'h00;
ROM_MEM[3561] <= 8'h97;
ROM_MEM[3562] <= 8'h45;
ROM_MEM[3563] <= 8'hFC;
ROM_MEM[3564] <= 8'h50;
ROM_MEM[3565] <= 8'h00;
ROM_MEM[3566] <= 8'h10;
ROM_MEM[3567] <= 8'h83;
ROM_MEM[3568] <= 8'h00;
ROM_MEM[3569] <= 8'h01;
ROM_MEM[3570] <= 8'h2D;
ROM_MEM[3571] <= 8'h6B;
ROM_MEM[3572] <= 8'hFD;
ROM_MEM[3573] <= 8'h47;
ROM_MEM[3574] <= 8'h04;
ROM_MEM[3575] <= 8'hFD;
ROM_MEM[3576] <= 8'h50;
ROM_MEM[3577] <= 8'h18;
ROM_MEM[3578] <= 8'hFC;
ROM_MEM[3579] <= 8'h50;
ROM_MEM[3580] <= 8'h02;
ROM_MEM[3581] <= 8'h2A;
ROM_MEM[3582] <= 8'h04;
ROM_MEM[3583] <= 8'h43;
ROM_MEM[3584] <= 8'h50;
ROM_MEM[3585] <= 8'h82;
ROM_MEM[3586] <= 8'hFF;
ROM_MEM[3587] <= 8'hB3;
ROM_MEM[3588] <= 8'h50;
ROM_MEM[3589] <= 8'h00;
ROM_MEM[3590] <= 8'h2C;
ROM_MEM[3591] <= 8'h57;
ROM_MEM[3592] <= 8'hFC;
ROM_MEM[3593] <= 8'h50;
ROM_MEM[3594] <= 8'h04;
ROM_MEM[3595] <= 8'h2A;
ROM_MEM[3596] <= 8'h04;
ROM_MEM[3597] <= 8'h43;
ROM_MEM[3598] <= 8'h50;
ROM_MEM[3599] <= 8'h82;
ROM_MEM[3600] <= 8'hFF;
ROM_MEM[3601] <= 8'hB3;
ROM_MEM[3602] <= 8'h50;
ROM_MEM[3603] <= 8'h00;
ROM_MEM[3604] <= 8'h2C;
ROM_MEM[3605] <= 8'h49;
ROM_MEM[3606] <= 8'hFC;
ROM_MEM[3607] <= 8'h47;
ROM_MEM[3608] <= 8'h00;
ROM_MEM[3609] <= 8'hFD;
ROM_MEM[3610] <= 8'h50;
ROM_MEM[3611] <= 8'h00;
ROM_MEM[3612] <= 8'h86;
ROM_MEM[3613] <= 8'h86;
ROM_MEM[3614] <= 8'hBD;
ROM_MEM[3615] <= 8'hCD;
ROM_MEM[3616] <= 8'hBA;
ROM_MEM[3617] <= 8'hFC;
ROM_MEM[3618] <= 8'h50;
ROM_MEM[3619] <= 8'h04;
ROM_MEM[3620] <= 8'hC3;
ROM_MEM[3621] <= 8'hFF;
ROM_MEM[3622] <= 8'h98;
ROM_MEM[3623] <= 8'h84;
ROM_MEM[3624] <= 8'h1F;
ROM_MEM[3625] <= 8'hED;
ROM_MEM[3626] <= 8'hA1;
ROM_MEM[3627] <= 8'hFC;
ROM_MEM[3628] <= 8'h50;
ROM_MEM[3629] <= 8'h02;
ROM_MEM[3630] <= 8'h84;
ROM_MEM[3631] <= 8'h1F;
ROM_MEM[3632] <= 8'hED;
ROM_MEM[3633] <= 8'hA1;
ROM_MEM[3634] <= 8'hCC;
ROM_MEM[3635] <= 8'h63;
ROM_MEM[3636] <= 8'hFF;
ROM_MEM[3637] <= 8'hED;
ROM_MEM[3638] <= 8'hA1;
ROM_MEM[3639] <= 8'h86;
ROM_MEM[3640] <= 8'h06;
ROM_MEM[3641] <= 8'h97;
ROM_MEM[3642] <= 8'h01;
ROM_MEM[3643] <= 8'hFC;
ROM_MEM[3644] <= 8'h50;
ROM_MEM[3645] <= 8'h18;
ROM_MEM[3646] <= 8'h0A;
ROM_MEM[3647] <= 8'h01;
ROM_MEM[3648] <= 8'h27;
ROM_MEM[3649] <= 8'h06;
ROM_MEM[3650] <= 8'h58;
ROM_MEM[3651] <= 8'h49;
ROM_MEM[3652] <= 8'h2A;
ROM_MEM[3653] <= 8'hF8;
ROM_MEM[3654] <= 8'h84;
ROM_MEM[3655] <= 8'h7F;
ROM_MEM[3656] <= 8'hD6;
ROM_MEM[3657] <= 8'h01;
ROM_MEM[3658] <= 8'hCA;
ROM_MEM[3659] <= 8'h70;
ROM_MEM[3660] <= 8'hE7;
ROM_MEM[3661] <= 8'hA0;
ROM_MEM[3662] <= 8'hA7;
ROM_MEM[3663] <= 8'hA0;
ROM_MEM[3664] <= 8'hCC;
ROM_MEM[3665] <= 8'hA0;
ROM_MEM[3666] <= 8'h16;
ROM_MEM[3667] <= 8'hED;
ROM_MEM[3668] <= 8'hA1;
ROM_MEM[3669] <= 8'hCC;
ROM_MEM[3670] <= 8'h72;
ROM_MEM[3671] <= 8'h00;
ROM_MEM[3672] <= 8'hED;
ROM_MEM[3673] <= 8'hA1;
ROM_MEM[3674] <= 8'hCC;
ROM_MEM[3675] <= 8'h80;
ROM_MEM[3676] <= 8'h40;
ROM_MEM[3677] <= 8'hED;
ROM_MEM[3678] <= 8'hA1;
ROM_MEM[3679] <= 8'h39;
ROM_MEM[3680] <= 8'h96;
ROM_MEM[3681] <= 8'hBD;
ROM_MEM[3682] <= 8'h2F;
ROM_MEM[3683] <= 8'h0A;
ROM_MEM[3684] <= 8'h0A;
ROM_MEM[3685] <= 8'hBD;
ROM_MEM[3686] <= 8'h86;
ROM_MEM[3687] <= 8'h00;
ROM_MEM[3688] <= 8'h97;
ROM_MEM[3689] <= 8'hB7;
ROM_MEM[3690] <= 8'h97;
ROM_MEM[3691] <= 8'hBC;
ROM_MEM[3692] <= 8'h20;
ROM_MEM[3693] <= 8'h04;
ROM_MEM[3694] <= 8'h86;
ROM_MEM[3695] <= 8'h00;
ROM_MEM[3696] <= 8'h97;
ROM_MEM[3697] <= 8'hBD;
ROM_MEM[3698] <= 8'h86;
ROM_MEM[3699] <= 8'h00;
ROM_MEM[3700] <= 8'h97;
ROM_MEM[3701] <= 8'hBC;
ROM_MEM[3702] <= 8'h1A;
ROM_MEM[3703] <= 8'h10;
ROM_MEM[3704] <= 8'h96;
ROM_MEM[3705] <= 8'h31;
ROM_MEM[3706] <= 8'h27;
ROM_MEM[3707] <= 8'h0B;
ROM_MEM[3708] <= 8'h7C;
ROM_MEM[3709] <= 8'h4B;
ROM_MEM[3710] <= 8'h1B;
ROM_MEM[3711] <= 8'h0F;
ROM_MEM[3712] <= 8'hBD;
ROM_MEM[3713] <= 8'hC6;
ROM_MEM[3714] <= 8'h08;
ROM_MEM[3715] <= 8'hD7;
ROM_MEM[3716] <= 8'hB7;
ROM_MEM[3717] <= 8'h0F;
ROM_MEM[3718] <= 8'h31;
ROM_MEM[3719] <= 8'h96;
ROM_MEM[3720] <= 8'hB7;
ROM_MEM[3721] <= 8'h2F;
ROM_MEM[3722] <= 8'h14;
ROM_MEM[3723] <= 8'h0A;
ROM_MEM[3724] <= 8'hB7;
ROM_MEM[3725] <= 8'h97;
ROM_MEM[3726] <= 8'hBC;
ROM_MEM[3727] <= 8'hDC;
ROM_MEM[3728] <= 8'h74;
ROM_MEM[3729] <= 8'hDD;
ROM_MEM[3730] <= 8'hB8;
ROM_MEM[3731] <= 8'hDC;
ROM_MEM[3732] <= 8'h6B;
ROM_MEM[3733] <= 8'hDD;
ROM_MEM[3734] <= 8'hBA;
ROM_MEM[3735] <= 8'hDC;
ROM_MEM[3736] <= 8'h2D;
ROM_MEM[3737] <= 8'hDD;
ROM_MEM[3738] <= 8'hB3;
ROM_MEM[3739] <= 8'hDC;
ROM_MEM[3740] <= 8'h2F;
ROM_MEM[3741] <= 8'hDD;
ROM_MEM[3742] <= 8'hB5;
ROM_MEM[3743] <= 8'h1C;
ROM_MEM[3744] <= 8'hEF;
ROM_MEM[3745] <= 8'h96;
ROM_MEM[3746] <= 8'hB7;
ROM_MEM[3747] <= 8'h81;
ROM_MEM[3748] <= 8'h07;
ROM_MEM[3749] <= 8'h26;
ROM_MEM[3750] <= 8'h0B;
ROM_MEM[3751] <= 8'hB6;
ROM_MEM[3752] <= 8'h4B;
ROM_MEM[3753] <= 8'h36;
ROM_MEM[3754] <= 8'h26;
ROM_MEM[3755] <= 8'h03;
ROM_MEM[3756] <= 8'h7A;
ROM_MEM[3757] <= 8'h4B;
ROM_MEM[3758] <= 8'h36;
ROM_MEM[3759] <= 8'hBD;
ROM_MEM[3760] <= 8'hBE;
ROM_MEM[3761] <= 8'h16;
ROM_MEM[3762] <= 8'h86;
ROM_MEM[3763] <= 8'hFF;
ROM_MEM[3764] <= 8'h97;
ROM_MEM[3765] <= 8'hC4;
ROM_MEM[3766] <= 8'h97;
ROM_MEM[3767] <= 8'hC8;
ROM_MEM[3768] <= 8'h97;
ROM_MEM[3769] <= 8'hCC;
ROM_MEM[3770] <= 8'h97;
ROM_MEM[3771] <= 8'hD0;
ROM_MEM[3772] <= 8'h39;
ROM_MEM[3773] <= 8'h96;
ROM_MEM[3774] <= 8'hBC;
ROM_MEM[3775] <= 8'h9A;
ROM_MEM[3776] <= 8'hBD;
ROM_MEM[3777] <= 8'h26;
ROM_MEM[3778] <= 8'h01;
ROM_MEM[3779] <= 8'h39;
ROM_MEM[3780] <= 8'hB6;
ROM_MEM[3781] <= 8'h4B;
ROM_MEM[3782] <= 8'h1B;
ROM_MEM[3783] <= 8'h84;
ROM_MEM[3784] <= 8'h01;
ROM_MEM[3785] <= 8'h27;
ROM_MEM[3786] <= 8'h5A;
ROM_MEM[3787] <= 8'hCC;
ROM_MEM[3788] <= 8'hFF;
ROM_MEM[3789] <= 8'h98;
ROM_MEM[3790] <= 8'hF3;
ROM_MEM[3791] <= 8'h4B;
ROM_MEM[3792] <= 8'h1E;
ROM_MEM[3793] <= 8'h84;
ROM_MEM[3794] <= 8'h1F;
ROM_MEM[3795] <= 8'hED;
ROM_MEM[3796] <= 8'hA1;
ROM_MEM[3797] <= 8'hDC;
ROM_MEM[3798] <= 8'hB5;
ROM_MEM[3799] <= 8'h83;
ROM_MEM[3800] <= 8'h00;
ROM_MEM[3801] <= 8'h00;
ROM_MEM[3802] <= 8'hB3;
ROM_MEM[3803] <= 8'h4B;
ROM_MEM[3804] <= 8'h1E;
ROM_MEM[3805] <= 8'hDD;
ROM_MEM[3806] <= 8'h03;
ROM_MEM[3807] <= 8'hCC;
ROM_MEM[3808] <= 8'hFE;
ROM_MEM[3809] <= 8'h7A;
ROM_MEM[3810] <= 8'hF3;
ROM_MEM[3811] <= 8'h4B;
ROM_MEM[3812] <= 8'h1C;
ROM_MEM[3813] <= 8'h84;
ROM_MEM[3814] <= 8'h1F;
ROM_MEM[3815] <= 8'hED;
ROM_MEM[3816] <= 8'hA1;
ROM_MEM[3817] <= 8'hDC;
ROM_MEM[3818] <= 8'hB3;
ROM_MEM[3819] <= 8'h83;
ROM_MEM[3820] <= 8'hFE;
ROM_MEM[3821] <= 8'h7A;
ROM_MEM[3822] <= 8'hB3;
ROM_MEM[3823] <= 8'h4B;
ROM_MEM[3824] <= 8'h1C;
ROM_MEM[3825] <= 8'hDD;
ROM_MEM[3826] <= 8'h01;
ROM_MEM[3827] <= 8'hC6;
ROM_MEM[3828] <= 8'h00;
ROM_MEM[3829] <= 8'hBD;
ROM_MEM[3830] <= 8'hAF;
ROM_MEM[3831] <= 8'h87;
ROM_MEM[3832] <= 8'hCC;
ROM_MEM[3833] <= 8'hFD;
ROM_MEM[3834] <= 8'hFB;
ROM_MEM[3835] <= 8'hF3;
ROM_MEM[3836] <= 8'h4B;
ROM_MEM[3837] <= 8'h1E;
ROM_MEM[3838] <= 8'h84;
ROM_MEM[3839] <= 8'h1F;
ROM_MEM[3840] <= 8'hED;
ROM_MEM[3841] <= 8'hA1;
ROM_MEM[3842] <= 8'hDC;
ROM_MEM[3843] <= 8'hB5;
ROM_MEM[3844] <= 8'h83;
ROM_MEM[3845] <= 8'hFE;
ROM_MEM[3846] <= 8'h63;
ROM_MEM[3847] <= 8'hB3;
ROM_MEM[3848] <= 8'h4B;
ROM_MEM[3849] <= 8'h1E;
ROM_MEM[3850] <= 8'hDD;
ROM_MEM[3851] <= 8'h03;
ROM_MEM[3852] <= 8'hCC;
ROM_MEM[3853] <= 8'hFE;
ROM_MEM[3854] <= 8'h75;
ROM_MEM[3855] <= 8'hF3;
ROM_MEM[3856] <= 8'h4B;
ROM_MEM[3857] <= 8'h1C;
ROM_MEM[3858] <= 8'h84;
ROM_MEM[3859] <= 8'h1F;
ROM_MEM[3860] <= 8'hED;
ROM_MEM[3861] <= 8'hA1;
ROM_MEM[3862] <= 8'hDC;
ROM_MEM[3863] <= 8'hB3;
ROM_MEM[3864] <= 8'h83;
ROM_MEM[3865] <= 8'hFE;
ROM_MEM[3866] <= 8'h75;
ROM_MEM[3867] <= 8'hB3;
ROM_MEM[3868] <= 8'h4B;
ROM_MEM[3869] <= 8'h1C;
ROM_MEM[3870] <= 8'hDD;
ROM_MEM[3871] <= 8'h01;
ROM_MEM[3872] <= 8'hC6;
ROM_MEM[3873] <= 8'h08;
ROM_MEM[3874] <= 8'hBD;
ROM_MEM[3875] <= 8'hAF;
ROM_MEM[3876] <= 8'h87;
ROM_MEM[3877] <= 8'hB6;
ROM_MEM[3878] <= 8'h4B;
ROM_MEM[3879] <= 8'h1B;
ROM_MEM[3880] <= 8'h84;
ROM_MEM[3881] <= 8'h01;
ROM_MEM[3882] <= 8'h26;
ROM_MEM[3883] <= 8'h5A;
ROM_MEM[3884] <= 8'hCC;
ROM_MEM[3885] <= 8'hFD;
ROM_MEM[3886] <= 8'hFB;
ROM_MEM[3887] <= 8'hF3;
ROM_MEM[3888] <= 8'h4B;
ROM_MEM[3889] <= 8'h1E;
ROM_MEM[3890] <= 8'h84;
ROM_MEM[3891] <= 8'h1F;
ROM_MEM[3892] <= 8'hED;
ROM_MEM[3893] <= 8'hA1;
ROM_MEM[3894] <= 8'hDC;
ROM_MEM[3895] <= 8'hB5;
ROM_MEM[3896] <= 8'h83;
ROM_MEM[3897] <= 8'hFE;
ROM_MEM[3898] <= 8'h63;
ROM_MEM[3899] <= 8'hB3;
ROM_MEM[3900] <= 8'h4B;
ROM_MEM[3901] <= 8'h1E;
ROM_MEM[3902] <= 8'hDD;
ROM_MEM[3903] <= 8'h03;
ROM_MEM[3904] <= 8'hCC;
ROM_MEM[3905] <= 8'h01;
ROM_MEM[3906] <= 8'h8B;
ROM_MEM[3907] <= 8'hF3;
ROM_MEM[3908] <= 8'h4B;
ROM_MEM[3909] <= 8'h1C;
ROM_MEM[3910] <= 8'h84;
ROM_MEM[3911] <= 8'h1F;
ROM_MEM[3912] <= 8'hED;
ROM_MEM[3913] <= 8'hA1;
ROM_MEM[3914] <= 8'hDC;
ROM_MEM[3915] <= 8'hB3;
ROM_MEM[3916] <= 8'h83;
ROM_MEM[3917] <= 8'h01;
ROM_MEM[3918] <= 8'h8B;
ROM_MEM[3919] <= 8'hB3;
ROM_MEM[3920] <= 8'h4B;
ROM_MEM[3921] <= 8'h1C;
ROM_MEM[3922] <= 8'hDD;
ROM_MEM[3923] <= 8'h01;
ROM_MEM[3924] <= 8'hC6;
ROM_MEM[3925] <= 8'h00;
ROM_MEM[3926] <= 8'hBD;
ROM_MEM[3927] <= 8'hAF;
ROM_MEM[3928] <= 8'h87;
ROM_MEM[3929] <= 8'hCC;
ROM_MEM[3930] <= 8'hFF;
ROM_MEM[3931] <= 8'h98;
ROM_MEM[3932] <= 8'hF3;
ROM_MEM[3933] <= 8'h4B;
ROM_MEM[3934] <= 8'h1E;
ROM_MEM[3935] <= 8'h84;
ROM_MEM[3936] <= 8'h1F;
ROM_MEM[3937] <= 8'hED;
ROM_MEM[3938] <= 8'hA1;
ROM_MEM[3939] <= 8'hDC;
ROM_MEM[3940] <= 8'hB5;
ROM_MEM[3941] <= 8'h83;
ROM_MEM[3942] <= 8'h00;
ROM_MEM[3943] <= 8'h00;
ROM_MEM[3944] <= 8'hB3;
ROM_MEM[3945] <= 8'h4B;
ROM_MEM[3946] <= 8'h1E;
ROM_MEM[3947] <= 8'hDD;
ROM_MEM[3948] <= 8'h03;
ROM_MEM[3949] <= 8'hCC;
ROM_MEM[3950] <= 8'h01;
ROM_MEM[3951] <= 8'h86;
ROM_MEM[3952] <= 8'hF3;
ROM_MEM[3953] <= 8'h4B;
ROM_MEM[3954] <= 8'h1C;
ROM_MEM[3955] <= 8'h84;
ROM_MEM[3956] <= 8'h1F;
ROM_MEM[3957] <= 8'hED;
ROM_MEM[3958] <= 8'hA1;
ROM_MEM[3959] <= 8'hDC;
ROM_MEM[3960] <= 8'hB3;
ROM_MEM[3961] <= 8'h83;
ROM_MEM[3962] <= 8'h01;
ROM_MEM[3963] <= 8'h86;
ROM_MEM[3964] <= 8'hB3;
ROM_MEM[3965] <= 8'h4B;
ROM_MEM[3966] <= 8'h1C;
ROM_MEM[3967] <= 8'hDD;
ROM_MEM[3968] <= 8'h01;
ROM_MEM[3969] <= 8'hC6;
ROM_MEM[3970] <= 8'h08;
ROM_MEM[3971] <= 8'hBD;
ROM_MEM[3972] <= 8'hAF;
ROM_MEM[3973] <= 8'h87;
ROM_MEM[3974] <= 8'h39;
ROM_MEM[3975] <= 8'hCE;
ROM_MEM[3976] <= 8'hB0;
ROM_MEM[3977] <= 8'h4F;
ROM_MEM[3978] <= 8'h33;
ROM_MEM[3979] <= 8'hC5;
ROM_MEM[3980] <= 8'h96;
ROM_MEM[3981] <= 8'hBD;
ROM_MEM[3982] <= 8'h2F;
ROM_MEM[3983] <= 8'h0A;
ROM_MEM[3984] <= 8'hC6;
ROM_MEM[3985] <= 8'h3F;
ROM_MEM[3986] <= 8'h3D;
ROM_MEM[3987] <= 8'h86;
ROM_MEM[3988] <= 8'h63;
ROM_MEM[3989] <= 8'hED;
ROM_MEM[3990] <= 8'hA1;
ROM_MEM[3991] <= 8'h7E;
ROM_MEM[3992] <= 8'hAF;
ROM_MEM[3993] <= 8'hEF;
ROM_MEM[3994] <= 8'h8E;
ROM_MEM[3995] <= 8'h4C;
ROM_MEM[3996] <= 8'h00;
ROM_MEM[3997] <= 8'hEC;
ROM_MEM[3998] <= 8'hC1;
ROM_MEM[3999] <= 8'hED;
ROM_MEM[4000] <= 8'hA1;
ROM_MEM[4001] <= 8'hDC;
ROM_MEM[4002] <= 8'h03;
ROM_MEM[4003] <= 8'h2B;
ROM_MEM[4004] <= 8'h03;
ROM_MEM[4005] <= 8'hC3;
ROM_MEM[4006] <= 8'h00;
ROM_MEM[4007] <= 8'h01;
ROM_MEM[4008] <= 8'h47;
ROM_MEM[4009] <= 8'h56;
ROM_MEM[4010] <= 8'hED;
ROM_MEM[4011] <= 8'hA4;
ROM_MEM[4012] <= 8'h43;
ROM_MEM[4013] <= 8'h50;
ROM_MEM[4014] <= 8'h82;
ROM_MEM[4015] <= 8'hFF;
ROM_MEM[4016] <= 8'hD3;
ROM_MEM[4017] <= 8'h03;
ROM_MEM[4018] <= 8'hDD;
ROM_MEM[4019] <= 8'h03;
ROM_MEM[4020] <= 8'hEC;
ROM_MEM[4021] <= 8'hA4;
ROM_MEM[4022] <= 8'h84;
ROM_MEM[4023] <= 8'h1F;
ROM_MEM[4024] <= 8'hED;
ROM_MEM[4025] <= 8'hA1;
ROM_MEM[4026] <= 8'hDC;
ROM_MEM[4027] <= 8'h01;
ROM_MEM[4028] <= 8'h2B;
ROM_MEM[4029] <= 8'h03;
ROM_MEM[4030] <= 8'hC3;
ROM_MEM[4031] <= 8'h00;
ROM_MEM[4032] <= 8'h01;
ROM_MEM[4033] <= 8'h47;
ROM_MEM[4034] <= 8'h56;
ROM_MEM[4035] <= 8'hED;
ROM_MEM[4036] <= 8'hA4;
ROM_MEM[4037] <= 8'h43;
ROM_MEM[4038] <= 8'h50;
ROM_MEM[4039] <= 8'h82;
ROM_MEM[4040] <= 8'hFF;
ROM_MEM[4041] <= 8'hD3;
ROM_MEM[4042] <= 8'h01;
ROM_MEM[4043] <= 8'hDD;
ROM_MEM[4044] <= 8'h01;
ROM_MEM[4045] <= 8'hEC;
ROM_MEM[4046] <= 8'hA4;
ROM_MEM[4047] <= 8'h8A;
ROM_MEM[4048] <= 8'hE0;
ROM_MEM[4049] <= 8'hED;
ROM_MEM[4050] <= 8'hA1;
ROM_MEM[4051] <= 8'hDC;
ROM_MEM[4052] <= 8'h01;
ROM_MEM[4053] <= 8'hC3;
ROM_MEM[4054] <= 8'h00;
ROM_MEM[4055] <= 8'h08;
ROM_MEM[4056] <= 8'h2D;
ROM_MEM[4057] <= 8'hC3;
ROM_MEM[4058] <= 8'h83;
ROM_MEM[4059] <= 8'h00;
ROM_MEM[4060] <= 8'h10;
ROM_MEM[4061] <= 8'h2E;
ROM_MEM[4062] <= 8'hBE;
ROM_MEM[4063] <= 8'hDC;
ROM_MEM[4064] <= 8'h03;
ROM_MEM[4065] <= 8'hC3;
ROM_MEM[4066] <= 8'h00;
ROM_MEM[4067] <= 8'h08;
ROM_MEM[4068] <= 8'h2D;
ROM_MEM[4069] <= 8'hB7;
ROM_MEM[4070] <= 8'h83;
ROM_MEM[4071] <= 8'h00;
ROM_MEM[4072] <= 8'h10;
ROM_MEM[4073] <= 8'h2E;
ROM_MEM[4074] <= 8'hB2;
ROM_MEM[4075] <= 8'hEC;
ROM_MEM[4076] <= 8'hC1;
ROM_MEM[4077] <= 8'hED;
ROM_MEM[4078] <= 8'hA1;
ROM_MEM[4079] <= 8'hDC;
ROM_MEM[4080] <= 8'h03;
ROM_MEM[4081] <= 8'h84;
ROM_MEM[4082] <= 8'h1F;
ROM_MEM[4083] <= 8'hED;
ROM_MEM[4084] <= 8'hA1;
ROM_MEM[4085] <= 8'hDC;
ROM_MEM[4086] <= 8'h01;
ROM_MEM[4087] <= 8'h8A;
ROM_MEM[4088] <= 8'hE0;
ROM_MEM[4089] <= 8'hED;
ROM_MEM[4090] <= 8'hA1;
ROM_MEM[4091] <= 8'h96;
ROM_MEM[4092] <= 8'hBD;
ROM_MEM[4093] <= 8'h2F;
ROM_MEM[4094] <= 8'h07;
ROM_MEM[4095] <= 8'hCC;
ROM_MEM[4096] <= 8'hA0;
ROM_MEM[4097] <= 8'h11;
ROM_MEM[4098] <= 8'hED;
ROM_MEM[4099] <= 8'hA1;
ROM_MEM[4100] <= 8'h20;
ROM_MEM[4101] <= 8'h3E;
ROM_MEM[4102] <= 8'h2C;
ROM_MEM[4103] <= 8'h3C;
ROM_MEM[4104] <= 8'hF6;
ROM_MEM[4105] <= 8'h4B;
ROM_MEM[4106] <= 8'h22;
ROM_MEM[4107] <= 8'h86;
ROM_MEM[4108] <= 8'h71;
ROM_MEM[4109] <= 8'hED;
ROM_MEM[4110] <= 8'hA1;
ROM_MEM[4111] <= 8'hFC;
ROM_MEM[4112] <= 8'h4B;
ROM_MEM[4113] <= 8'h20;
ROM_MEM[4114] <= 8'hED;
ROM_MEM[4115] <= 8'hA1;
ROM_MEM[4116] <= 8'hB6;
ROM_MEM[4117] <= 8'h4B;
ROM_MEM[4118] <= 8'h23;
ROM_MEM[4119] <= 8'h84;
ROM_MEM[4120] <= 8'h01;
ROM_MEM[4121] <= 8'h27;
ROM_MEM[4122] <= 8'h05;
ROM_MEM[4123] <= 8'hCC;
ROM_MEM[4124] <= 8'hA0;
ROM_MEM[4125] <= 8'h1C;
ROM_MEM[4126] <= 8'hED;
ROM_MEM[4127] <= 8'hA1;
ROM_MEM[4128] <= 8'hB6;
ROM_MEM[4129] <= 8'h4B;
ROM_MEM[4130] <= 8'h23;
ROM_MEM[4131] <= 8'h84;
ROM_MEM[4132] <= 8'h02;
ROM_MEM[4133] <= 8'h27;
ROM_MEM[4134] <= 8'h05;
ROM_MEM[4135] <= 8'hCC;
ROM_MEM[4136] <= 8'hA0;
ROM_MEM[4137] <= 8'h23;
ROM_MEM[4138] <= 8'hED;
ROM_MEM[4139] <= 8'hA1;
ROM_MEM[4140] <= 8'hB6;
ROM_MEM[4141] <= 8'h4B;
ROM_MEM[4142] <= 8'h23;
ROM_MEM[4143] <= 8'h84;
ROM_MEM[4144] <= 8'h04;
ROM_MEM[4145] <= 8'h27;
ROM_MEM[4146] <= 8'h05;
ROM_MEM[4147] <= 8'hCC;
ROM_MEM[4148] <= 8'hA0;
ROM_MEM[4149] <= 8'h2A;
ROM_MEM[4150] <= 8'hED;
ROM_MEM[4151] <= 8'hA1;
ROM_MEM[4152] <= 8'hB6;
ROM_MEM[4153] <= 8'h4B;
ROM_MEM[4154] <= 8'h23;
ROM_MEM[4155] <= 8'h84;
ROM_MEM[4156] <= 8'h08;
ROM_MEM[4157] <= 8'h27;
ROM_MEM[4158] <= 8'h05;
ROM_MEM[4159] <= 8'hCC;
ROM_MEM[4160] <= 8'hA0;
ROM_MEM[4161] <= 8'h31;
ROM_MEM[4162] <= 8'hED;
ROM_MEM[4163] <= 8'hA1;
ROM_MEM[4164] <= 8'hCC;
ROM_MEM[4165] <= 8'h72;
ROM_MEM[4166] <= 8'h00;
ROM_MEM[4167] <= 8'hED;
ROM_MEM[4168] <= 8'hA1;
ROM_MEM[4169] <= 8'hCC;
ROM_MEM[4170] <= 8'h80;
ROM_MEM[4171] <= 8'h40;
ROM_MEM[4172] <= 8'hED;
ROM_MEM[4173] <= 8'hA1;
ROM_MEM[4174] <= 8'h39;
ROM_MEM[4175] <= 8'hA0;
ROM_MEM[4176] <= 8'h01;
ROM_MEM[4177] <= 8'hA0;
ROM_MEM[4178] <= 8'h02;
ROM_MEM[4179] <= 8'hA0;
ROM_MEM[4180] <= 8'h03;
ROM_MEM[4181] <= 8'hA0;
ROM_MEM[4182] <= 8'h04;
ROM_MEM[4183] <= 8'hA0;
ROM_MEM[4184] <= 8'h05;
ROM_MEM[4185] <= 8'hA0;
ROM_MEM[4186] <= 8'h06;
ROM_MEM[4187] <= 8'hA0;
ROM_MEM[4188] <= 8'h07;
ROM_MEM[4189] <= 8'hA0;
ROM_MEM[4190] <= 8'h08;
ROM_MEM[4191] <= 8'hA0;
ROM_MEM[4192] <= 8'h09;
ROM_MEM[4193] <= 8'hA0;
ROM_MEM[4194] <= 8'h0A;
ROM_MEM[4195] <= 8'hA0;
ROM_MEM[4196] <= 8'h0B;
ROM_MEM[4197] <= 8'hA0;
ROM_MEM[4198] <= 8'h0C;
ROM_MEM[4199] <= 8'hA0;
ROM_MEM[4200] <= 8'h0D;
ROM_MEM[4201] <= 8'hA0;
ROM_MEM[4202] <= 8'h0E;
ROM_MEM[4203] <= 8'hA0;
ROM_MEM[4204] <= 8'h0F;
ROM_MEM[4205] <= 8'hA0;
ROM_MEM[4206] <= 8'h10;
ROM_MEM[4207] <= 8'hA0;
ROM_MEM[4208] <= 8'h01;
ROM_MEM[4209] <= 8'h96;
ROM_MEM[4210] <= 8'hBC;
ROM_MEM[4211] <= 8'h27;
ROM_MEM[4212] <= 8'h1F;
ROM_MEM[4213] <= 8'hBD;
ROM_MEM[4214] <= 8'hB0;
ROM_MEM[4215] <= 8'h95;
ROM_MEM[4216] <= 8'hCC;
ROM_MEM[4217] <= 8'h02;
ROM_MEM[4218] <= 8'h00;
ROM_MEM[4219] <= 8'hFD;
ROM_MEM[4220] <= 8'h47;
ROM_MEM[4221] <= 8'h06;
ROM_MEM[4222] <= 8'hDC;
ROM_MEM[4223] <= 8'hCC;
ROM_MEM[4224] <= 8'h2B;
ROM_MEM[4225] <= 8'h07;
ROM_MEM[4226] <= 8'h86;
ROM_MEM[4227] <= 8'h04;
ROM_MEM[4228] <= 8'h97;
ROM_MEM[4229] <= 8'hBD;
ROM_MEM[4230] <= 8'hBD;
ROM_MEM[4231] <= 8'hAD;
ROM_MEM[4232] <= 8'h20;
ROM_MEM[4233] <= 8'h96;
ROM_MEM[4234] <= 8'h44;
ROM_MEM[4235] <= 8'h2F;
ROM_MEM[4236] <= 8'h07;
ROM_MEM[4237] <= 8'h86;
ROM_MEM[4238] <= 8'hFF;
ROM_MEM[4239] <= 8'h97;
ROM_MEM[4240] <= 8'h44;
ROM_MEM[4241] <= 8'hBD;
ROM_MEM[4242] <= 8'hAD;
ROM_MEM[4243] <= 8'h3E;
ROM_MEM[4244] <= 8'h39;
ROM_MEM[4245] <= 8'hCC;
ROM_MEM[4246] <= 8'h70;
ROM_MEM[4247] <= 8'h00;
ROM_MEM[4248] <= 8'hF3;
ROM_MEM[4249] <= 8'h50;
ROM_MEM[4250] <= 8'h40;
ROM_MEM[4251] <= 8'hDD;
ROM_MEM[4252] <= 8'h01;
ROM_MEM[4253] <= 8'hCC;
ROM_MEM[4254] <= 8'h00;
ROM_MEM[4255] <= 8'h00;
ROM_MEM[4256] <= 8'h93;
ROM_MEM[4257] <= 8'hB8;
ROM_MEM[4258] <= 8'hBD;
ROM_MEM[4259] <= 8'hCD;
ROM_MEM[4260] <= 8'hA2;
ROM_MEM[4261] <= 8'hD3;
ROM_MEM[4262] <= 8'hB8;
ROM_MEM[4263] <= 8'hF3;
ROM_MEM[4264] <= 8'h50;
ROM_MEM[4265] <= 8'h42;
ROM_MEM[4266] <= 8'hDD;
ROM_MEM[4267] <= 8'h03;
ROM_MEM[4268] <= 8'hCC;
ROM_MEM[4269] <= 8'h00;
ROM_MEM[4270] <= 8'h00;
ROM_MEM[4271] <= 8'h93;
ROM_MEM[4272] <= 8'hBA;
ROM_MEM[4273] <= 8'hBD;
ROM_MEM[4274] <= 8'hCD;
ROM_MEM[4275] <= 8'hA2;
ROM_MEM[4276] <= 8'hD3;
ROM_MEM[4277] <= 8'hBA;
ROM_MEM[4278] <= 8'hF3;
ROM_MEM[4279] <= 8'h50;
ROM_MEM[4280] <= 8'h44;
ROM_MEM[4281] <= 8'hDD;
ROM_MEM[4282] <= 8'h05;
ROM_MEM[4283] <= 8'hCC;
ROM_MEM[4284] <= 8'hF0;
ROM_MEM[4285] <= 8'h00;
ROM_MEM[4286] <= 8'h93;
ROM_MEM[4287] <= 8'h05;
ROM_MEM[4288] <= 8'h10;
ROM_MEM[4289] <= 8'h2D;
ROM_MEM[4290] <= 8'h00;
ROM_MEM[4291] <= 8'h94;
ROM_MEM[4292] <= 8'hFD;
ROM_MEM[4293] <= 8'h47;
ROM_MEM[4294] <= 8'h06;
ROM_MEM[4295] <= 8'hFC;
ROM_MEM[4296] <= 8'h50;
ROM_MEM[4297] <= 8'h44;
ROM_MEM[4298] <= 8'h93;
ROM_MEM[4299] <= 8'h05;
ROM_MEM[4300] <= 8'hFD;
ROM_MEM[4301] <= 8'h47;
ROM_MEM[4302] <= 8'h04;
ROM_MEM[4303] <= 8'hDC;
ROM_MEM[4304] <= 8'h03;
ROM_MEM[4305] <= 8'hB3;
ROM_MEM[4306] <= 8'h50;
ROM_MEM[4307] <= 8'h42;
ROM_MEM[4308] <= 8'hFD;
ROM_MEM[4309] <= 8'h50;
ROM_MEM[4310] <= 8'h02;
ROM_MEM[4311] <= 8'hDC;
ROM_MEM[4312] <= 8'h01;
ROM_MEM[4313] <= 8'hB3;
ROM_MEM[4314] <= 8'h50;
ROM_MEM[4315] <= 8'h40;
ROM_MEM[4316] <= 8'hFD;
ROM_MEM[4317] <= 8'h50;
ROM_MEM[4318] <= 8'h04;
ROM_MEM[4319] <= 8'hFC;
ROM_MEM[4320] <= 8'h47;
ROM_MEM[4321] <= 8'h00;
ROM_MEM[4322] <= 8'hFD;
ROM_MEM[4323] <= 8'h50;
ROM_MEM[4324] <= 8'h00;
ROM_MEM[4325] <= 8'h86;
ROM_MEM[4326] <= 8'h86;
ROM_MEM[4327] <= 8'hBD;
ROM_MEM[4328] <= 8'hCD;
ROM_MEM[4329] <= 8'hBA;
ROM_MEM[4330] <= 8'hDC;
ROM_MEM[4331] <= 8'h03;
ROM_MEM[4332] <= 8'hB3;
ROM_MEM[4333] <= 8'h50;
ROM_MEM[4334] <= 8'h02;
ROM_MEM[4335] <= 8'h2B;
ROM_MEM[4336] <= 8'h08;
ROM_MEM[4337] <= 8'h10;
ROM_MEM[4338] <= 8'h83;
ROM_MEM[4339] <= 8'h04;
ROM_MEM[4340] <= 8'h00;
ROM_MEM[4341] <= 8'h2E;
ROM_MEM[4342] <= 8'h61;
ROM_MEM[4343] <= 8'h20;
ROM_MEM[4344] <= 8'h06;
ROM_MEM[4345] <= 8'h10;
ROM_MEM[4346] <= 8'h83;
ROM_MEM[4347] <= 8'hFC;
ROM_MEM[4348] <= 8'h00;
ROM_MEM[4349] <= 8'h2D;
ROM_MEM[4350] <= 8'h59;
ROM_MEM[4351] <= 8'hDD;
ROM_MEM[4352] <= 8'h03;
ROM_MEM[4353] <= 8'hDC;
ROM_MEM[4354] <= 8'h01;
ROM_MEM[4355] <= 8'hB3;
ROM_MEM[4356] <= 8'h50;
ROM_MEM[4357] <= 8'h04;
ROM_MEM[4358] <= 8'hDD;
ROM_MEM[4359] <= 8'h01;
ROM_MEM[4360] <= 8'hDD;
ROM_MEM[4361] <= 8'hC0;
ROM_MEM[4362] <= 8'hCC;
ROM_MEM[4363] <= 8'hF0;
ROM_MEM[4364] <= 8'h00;
ROM_MEM[4365] <= 8'hDD;
ROM_MEM[4366] <= 8'h05;
ROM_MEM[4367] <= 8'h86;
ROM_MEM[4368] <= 8'hFF;
ROM_MEM[4369] <= 8'h97;
ROM_MEM[4370] <= 8'hBD;
ROM_MEM[4371] <= 8'h86;
ROM_MEM[4372] <= 8'h03;
ROM_MEM[4373] <= 8'hB7;
ROM_MEM[4374] <= 8'h4B;
ROM_MEM[4375] <= 8'h23;
ROM_MEM[4376] <= 8'h96;
ROM_MEM[4377] <= 8'h01;
ROM_MEM[4378] <= 8'hB0;
ROM_MEM[4379] <= 8'h50;
ROM_MEM[4380] <= 8'h40;
ROM_MEM[4381] <= 8'hC6;
ROM_MEM[4382] <= 8'h03;
ROM_MEM[4383] <= 8'h3D;
ROM_MEM[4384] <= 8'h10;
ROM_MEM[4385] <= 8'h83;
ROM_MEM[4386] <= 8'h00;
ROM_MEM[4387] <= 8'hE0;
ROM_MEM[4388] <= 8'h25;
ROM_MEM[4389] <= 8'h02;
ROM_MEM[4390] <= 8'hC6;
ROM_MEM[4391] <= 8'hE0;
ROM_MEM[4392] <= 8'hF7;
ROM_MEM[4393] <= 8'h4B;
ROM_MEM[4394] <= 8'h22;
ROM_MEM[4395] <= 8'hCC;
ROM_MEM[4396] <= 8'h62;
ROM_MEM[4397] <= 8'h80;
ROM_MEM[4398] <= 8'hFD;
ROM_MEM[4399] <= 8'h4B;
ROM_MEM[4400] <= 8'h20;
ROM_MEM[4401] <= 8'h96;
ROM_MEM[4402] <= 8'h95;
ROM_MEM[4403] <= 8'h27;
ROM_MEM[4404] <= 8'h22;
ROM_MEM[4405] <= 8'h96;
ROM_MEM[4406] <= 8'h44;
ROM_MEM[4407] <= 8'h26;
ROM_MEM[4408] <= 8'h1E;
ROM_MEM[4409] <= 8'hDC;
ROM_MEM[4410] <= 8'h03;
ROM_MEM[4411] <= 8'hC3;
ROM_MEM[4412] <= 8'h02;
ROM_MEM[4413] <= 8'h00;
ROM_MEM[4414] <= 8'h2D;
ROM_MEM[4415] <= 8'h17;
ROM_MEM[4416] <= 8'h83;
ROM_MEM[4417] <= 8'h04;
ROM_MEM[4418] <= 8'h00;
ROM_MEM[4419] <= 8'h2E;
ROM_MEM[4420] <= 8'h12;
ROM_MEM[4421] <= 8'hDC;
ROM_MEM[4422] <= 8'h01;
ROM_MEM[4423] <= 8'h93;
ROM_MEM[4424] <= 8'h96;
ROM_MEM[4425] <= 8'hC3;
ROM_MEM[4426] <= 8'h02;
ROM_MEM[4427] <= 8'h00;
ROM_MEM[4428] <= 8'h2D;
ROM_MEM[4429] <= 8'h09;
ROM_MEM[4430] <= 8'h83;
ROM_MEM[4431] <= 8'h04;
ROM_MEM[4432] <= 8'h00;
ROM_MEM[4433] <= 8'h2E;
ROM_MEM[4434] <= 8'h04;
ROM_MEM[4435] <= 8'h86;
ROM_MEM[4436] <= 8'h01;
ROM_MEM[4437] <= 8'h97;
ROM_MEM[4438] <= 8'h44;
ROM_MEM[4439] <= 8'h39;
ROM_MEM[4440] <= 8'hDC;
ROM_MEM[4441] <= 8'h03;
ROM_MEM[4442] <= 8'h10;
ROM_MEM[4443] <= 8'h2A;
ROM_MEM[4444] <= 8'h00;
ROM_MEM[4445] <= 8'h85;
ROM_MEM[4446] <= 8'hCC;
ROM_MEM[4447] <= 8'hFC;
ROM_MEM[4448] <= 8'h00;
ROM_MEM[4449] <= 8'h93;
ROM_MEM[4450] <= 8'h03;
ROM_MEM[4451] <= 8'h10;
ROM_MEM[4452] <= 8'h2D;
ROM_MEM[4453] <= 8'h00;
ROM_MEM[4454] <= 8'hF9;
ROM_MEM[4455] <= 8'hFD;
ROM_MEM[4456] <= 8'h47;
ROM_MEM[4457] <= 8'h06;
ROM_MEM[4458] <= 8'hFC;
ROM_MEM[4459] <= 8'h50;
ROM_MEM[4460] <= 8'h42;
ROM_MEM[4461] <= 8'h93;
ROM_MEM[4462] <= 8'h03;
ROM_MEM[4463] <= 8'hFD;
ROM_MEM[4464] <= 8'h47;
ROM_MEM[4465] <= 8'h04;
ROM_MEM[4466] <= 8'hDC;
ROM_MEM[4467] <= 8'h05;
ROM_MEM[4468] <= 8'hB3;
ROM_MEM[4469] <= 8'h50;
ROM_MEM[4470] <= 8'h44;
ROM_MEM[4471] <= 8'hFD;
ROM_MEM[4472] <= 8'h50;
ROM_MEM[4473] <= 8'h04;
ROM_MEM[4474] <= 8'hDC;
ROM_MEM[4475] <= 8'h01;
ROM_MEM[4476] <= 8'hB3;
ROM_MEM[4477] <= 8'h50;
ROM_MEM[4478] <= 8'h40;
ROM_MEM[4479] <= 8'hFD;
ROM_MEM[4480] <= 8'h50;
ROM_MEM[4481] <= 8'h02;
ROM_MEM[4482] <= 8'hFC;
ROM_MEM[4483] <= 8'h47;
ROM_MEM[4484] <= 8'h00;
ROM_MEM[4485] <= 8'hFD;
ROM_MEM[4486] <= 8'h50;
ROM_MEM[4487] <= 8'h00;
ROM_MEM[4488] <= 8'h86;
ROM_MEM[4489] <= 8'h86;
ROM_MEM[4490] <= 8'hBD;
ROM_MEM[4491] <= 8'hCD;
ROM_MEM[4492] <= 8'hBA;
ROM_MEM[4493] <= 8'hDC;
ROM_MEM[4494] <= 8'h05;
ROM_MEM[4495] <= 8'hB3;
ROM_MEM[4496] <= 8'h50;
ROM_MEM[4497] <= 8'h04;
ROM_MEM[4498] <= 8'h2B;
ROM_MEM[4499] <= 8'h0A;
ROM_MEM[4500] <= 8'h10;
ROM_MEM[4501] <= 8'h83;
ROM_MEM[4502] <= 8'h00;
ROM_MEM[4503] <= 8'h00;
ROM_MEM[4504] <= 8'h10;
ROM_MEM[4505] <= 8'h2E;
ROM_MEM[4506] <= 8'h00;
ROM_MEM[4507] <= 8'hC4;
ROM_MEM[4508] <= 8'h20;
ROM_MEM[4509] <= 8'h08;
ROM_MEM[4510] <= 8'h10;
ROM_MEM[4511] <= 8'h83;
ROM_MEM[4512] <= 8'hF0;
ROM_MEM[4513] <= 8'h00;
ROM_MEM[4514] <= 8'h10;
ROM_MEM[4515] <= 8'h2D;
ROM_MEM[4516] <= 8'h00;
ROM_MEM[4517] <= 8'hBA;
ROM_MEM[4518] <= 8'hDD;
ROM_MEM[4519] <= 8'h05;
ROM_MEM[4520] <= 8'hC3;
ROM_MEM[4521] <= 8'h10;
ROM_MEM[4522] <= 8'h00;
ROM_MEM[4523] <= 8'hDD;
ROM_MEM[4524] <= 8'hBE;
ROM_MEM[4525] <= 8'hDC;
ROM_MEM[4526] <= 8'h01;
ROM_MEM[4527] <= 8'hB3;
ROM_MEM[4528] <= 8'h50;
ROM_MEM[4529] <= 8'h02;
ROM_MEM[4530] <= 8'hDD;
ROM_MEM[4531] <= 8'h01;
ROM_MEM[4532] <= 8'hDD;
ROM_MEM[4533] <= 8'hC0;
ROM_MEM[4534] <= 8'hCC;
ROM_MEM[4535] <= 8'hFC;
ROM_MEM[4536] <= 8'h00;
ROM_MEM[4537] <= 8'hDD;
ROM_MEM[4538] <= 8'h03;
ROM_MEM[4539] <= 8'h86;
ROM_MEM[4540] <= 8'hFF;
ROM_MEM[4541] <= 8'h97;
ROM_MEM[4542] <= 8'hBD;
ROM_MEM[4543] <= 8'h86;
ROM_MEM[4544] <= 8'h09;
ROM_MEM[4545] <= 8'hB7;
ROM_MEM[4546] <= 8'h4B;
ROM_MEM[4547] <= 8'h23;
ROM_MEM[4548] <= 8'h96;
ROM_MEM[4549] <= 8'h01;
ROM_MEM[4550] <= 8'hB0;
ROM_MEM[4551] <= 8'h50;
ROM_MEM[4552] <= 8'h40;
ROM_MEM[4553] <= 8'hC6;
ROM_MEM[4554] <= 8'h03;
ROM_MEM[4555] <= 8'h3D;
ROM_MEM[4556] <= 8'h10;
ROM_MEM[4557] <= 8'h83;
ROM_MEM[4558] <= 8'h00;
ROM_MEM[4559] <= 8'hE0;
ROM_MEM[4560] <= 8'h25;
ROM_MEM[4561] <= 8'h02;
ROM_MEM[4562] <= 8'hC6;
ROM_MEM[4563] <= 8'hE0;
ROM_MEM[4564] <= 8'hF7;
ROM_MEM[4565] <= 8'h4B;
ROM_MEM[4566] <= 8'h22;
ROM_MEM[4567] <= 8'hCC;
ROM_MEM[4568] <= 8'h62;
ROM_MEM[4569] <= 8'h80;
ROM_MEM[4570] <= 8'hFD;
ROM_MEM[4571] <= 8'h4B;
ROM_MEM[4572] <= 8'h20;
ROM_MEM[4573] <= 8'h8E;
ROM_MEM[4574] <= 8'h49;
ROM_MEM[4575] <= 8'h89;
ROM_MEM[4576] <= 8'h7E;
ROM_MEM[4577] <= 8'hB2;
ROM_MEM[4578] <= 8'h61;
ROM_MEM[4579] <= 8'h83;
ROM_MEM[4580] <= 8'h04;
ROM_MEM[4581] <= 8'h00;
ROM_MEM[4582] <= 8'h2D;
ROM_MEM[4583] <= 8'h78;
ROM_MEM[4584] <= 8'hFD;
ROM_MEM[4585] <= 8'h47;
ROM_MEM[4586] <= 8'h06;
ROM_MEM[4587] <= 8'hDC;
ROM_MEM[4588] <= 8'h03;
ROM_MEM[4589] <= 8'hB3;
ROM_MEM[4590] <= 8'h50;
ROM_MEM[4591] <= 8'h42;
ROM_MEM[4592] <= 8'hFD;
ROM_MEM[4593] <= 8'h47;
ROM_MEM[4594] <= 8'h04;
ROM_MEM[4595] <= 8'hDC;
ROM_MEM[4596] <= 8'h05;
ROM_MEM[4597] <= 8'hB3;
ROM_MEM[4598] <= 8'h50;
ROM_MEM[4599] <= 8'h44;
ROM_MEM[4600] <= 8'hFD;
ROM_MEM[4601] <= 8'h50;
ROM_MEM[4602] <= 8'h04;
ROM_MEM[4603] <= 8'hDC;
ROM_MEM[4604] <= 8'h01;
ROM_MEM[4605] <= 8'hB3;
ROM_MEM[4606] <= 8'h50;
ROM_MEM[4607] <= 8'h40;
ROM_MEM[4608] <= 8'hFD;
ROM_MEM[4609] <= 8'h50;
ROM_MEM[4610] <= 8'h02;
ROM_MEM[4611] <= 8'hFC;
ROM_MEM[4612] <= 8'h47;
ROM_MEM[4613] <= 8'h00;
ROM_MEM[4614] <= 8'hFD;
ROM_MEM[4615] <= 8'h50;
ROM_MEM[4616] <= 8'h00;
ROM_MEM[4617] <= 8'h86;
ROM_MEM[4618] <= 8'h86;
ROM_MEM[4619] <= 8'hBD;
ROM_MEM[4620] <= 8'hCD;
ROM_MEM[4621] <= 8'hBA;
ROM_MEM[4622] <= 8'hDC;
ROM_MEM[4623] <= 8'h05;
ROM_MEM[4624] <= 8'hB3;
ROM_MEM[4625] <= 8'h50;
ROM_MEM[4626] <= 8'h04;
ROM_MEM[4627] <= 8'h2B;
ROM_MEM[4628] <= 8'h08;
ROM_MEM[4629] <= 8'h10;
ROM_MEM[4630] <= 8'h83;
ROM_MEM[4631] <= 8'h00;
ROM_MEM[4632] <= 8'h00;
ROM_MEM[4633] <= 8'h2E;
ROM_MEM[4634] <= 8'h45;
ROM_MEM[4635] <= 8'h20;
ROM_MEM[4636] <= 8'h06;
ROM_MEM[4637] <= 8'h10;
ROM_MEM[4638] <= 8'h83;
ROM_MEM[4639] <= 8'hF0;
ROM_MEM[4640] <= 8'h00;
ROM_MEM[4641] <= 8'h2D;
ROM_MEM[4642] <= 8'h3D;
ROM_MEM[4643] <= 8'hDD;
ROM_MEM[4644] <= 8'h05;
ROM_MEM[4645] <= 8'hC3;
ROM_MEM[4646] <= 8'h10;
ROM_MEM[4647] <= 8'h00;
ROM_MEM[4648] <= 8'hDD;
ROM_MEM[4649] <= 8'hBE;
ROM_MEM[4650] <= 8'hDC;
ROM_MEM[4651] <= 8'h01;
ROM_MEM[4652] <= 8'hB3;
ROM_MEM[4653] <= 8'h50;
ROM_MEM[4654] <= 8'h02;
ROM_MEM[4655] <= 8'hDD;
ROM_MEM[4656] <= 8'h01;
ROM_MEM[4657] <= 8'hDD;
ROM_MEM[4658] <= 8'hC0;
ROM_MEM[4659] <= 8'hCC;
ROM_MEM[4660] <= 8'h04;
ROM_MEM[4661] <= 8'h00;
ROM_MEM[4662] <= 8'hDD;
ROM_MEM[4663] <= 8'h03;
ROM_MEM[4664] <= 8'h86;
ROM_MEM[4665] <= 8'hFF;
ROM_MEM[4666] <= 8'h97;
ROM_MEM[4667] <= 8'hBD;
ROM_MEM[4668] <= 8'h86;
ROM_MEM[4669] <= 8'h06;
ROM_MEM[4670] <= 8'hB7;
ROM_MEM[4671] <= 8'h4B;
ROM_MEM[4672] <= 8'h23;
ROM_MEM[4673] <= 8'h96;
ROM_MEM[4674] <= 8'h01;
ROM_MEM[4675] <= 8'hB0;
ROM_MEM[4676] <= 8'h50;
ROM_MEM[4677] <= 8'h40;
ROM_MEM[4678] <= 8'hC6;
ROM_MEM[4679] <= 8'h03;
ROM_MEM[4680] <= 8'h3D;
ROM_MEM[4681] <= 8'h10;
ROM_MEM[4682] <= 8'h83;
ROM_MEM[4683] <= 8'h00;
ROM_MEM[4684] <= 8'hE0;
ROM_MEM[4685] <= 8'h25;
ROM_MEM[4686] <= 8'h02;
ROM_MEM[4687] <= 8'hC6;
ROM_MEM[4688] <= 8'hE0;
ROM_MEM[4689] <= 8'hF7;
ROM_MEM[4690] <= 8'h4B;
ROM_MEM[4691] <= 8'h22;
ROM_MEM[4692] <= 8'hCC;
ROM_MEM[4693] <= 8'h62;
ROM_MEM[4694] <= 8'h80;
ROM_MEM[4695] <= 8'hFD;
ROM_MEM[4696] <= 8'h4B;
ROM_MEM[4697] <= 8'h20;
ROM_MEM[4698] <= 8'h8E;
ROM_MEM[4699] <= 8'h49;
ROM_MEM[4700] <= 8'h99;
ROM_MEM[4701] <= 8'h7E;
ROM_MEM[4702] <= 8'hB2;
ROM_MEM[4703] <= 8'h61;
ROM_MEM[4704] <= 8'h39;
ROM_MEM[4705] <= 8'h96;
ROM_MEM[4706] <= 8'hBC;
ROM_MEM[4707] <= 8'h26;
ROM_MEM[4708] <= 8'h01;
ROM_MEM[4709] <= 8'h39;
ROM_MEM[4710] <= 8'hD6;
ROM_MEM[4711] <= 8'hC0;
ROM_MEM[4712] <= 8'h54;
ROM_MEM[4713] <= 8'h54;
ROM_MEM[4714] <= 8'h54;
ROM_MEM[4715] <= 8'hC4;
ROM_MEM[4716] <= 8'h0F;
ROM_MEM[4717] <= 8'h3A;
ROM_MEM[4718] <= 8'hDC;
ROM_MEM[4719] <= 8'hC0;
ROM_MEM[4720] <= 8'h84;
ROM_MEM[4721] <= 8'h07;
ROM_MEM[4722] <= 8'h83;
ROM_MEM[4723] <= 8'h01;
ROM_MEM[4724] <= 8'hC0;
ROM_MEM[4725] <= 8'h2D;
ROM_MEM[4726] <= 8'h24;
ROM_MEM[4727] <= 8'h83;
ROM_MEM[4728] <= 8'h04;
ROM_MEM[4729] <= 8'h80;
ROM_MEM[4730] <= 8'h2E;
ROM_MEM[4731] <= 8'h1F;
ROM_MEM[4732] <= 8'h86;
ROM_MEM[4733] <= 8'h03;
ROM_MEM[4734] <= 8'h97;
ROM_MEM[4735] <= 8'h01;
ROM_MEM[4736] <= 8'hDC;
ROM_MEM[4737] <= 8'hBE;
ROM_MEM[4738] <= 8'h83;
ROM_MEM[4739] <= 8'h00;
ROM_MEM[4740] <= 8'h40;
ROM_MEM[4741] <= 8'h83;
ROM_MEM[4742] <= 8'h03;
ROM_MEM[4743] <= 8'h80;
ROM_MEM[4744] <= 8'h2E;
ROM_MEM[4745] <= 8'h08;
ROM_MEM[4746] <= 8'h83;
ROM_MEM[4747] <= 8'hFC;
ROM_MEM[4748] <= 8'h80;
ROM_MEM[4749] <= 8'h2D;
ROM_MEM[4750] <= 8'h0C;
ROM_MEM[4751] <= 8'h7E;
ROM_MEM[4752] <= 8'hB2;
ROM_MEM[4753] <= 8'h9C;
ROM_MEM[4754] <= 8'h83;
ROM_MEM[4755] <= 8'h00;
ROM_MEM[4756] <= 8'h80;
ROM_MEM[4757] <= 8'h08;
ROM_MEM[4758] <= 8'h01;
ROM_MEM[4759] <= 8'h08;
ROM_MEM[4760] <= 8'h01;
ROM_MEM[4761] <= 8'h26;
ROM_MEM[4762] <= 8'hEA;
ROM_MEM[4763] <= 8'h39;
ROM_MEM[4764] <= 8'h96;
ROM_MEM[4765] <= 8'h01;
ROM_MEM[4766] <= 8'hA4;
ROM_MEM[4767] <= 8'h84;
ROM_MEM[4768] <= 8'h27;
ROM_MEM[4769] <= 8'h2F;
ROM_MEM[4770] <= 8'h97;
ROM_MEM[4771] <= 8'h02;
ROM_MEM[4772] <= 8'h96;
ROM_MEM[4773] <= 8'h01;
ROM_MEM[4774] <= 8'h48;
ROM_MEM[4775] <= 8'h94;
ROM_MEM[4776] <= 8'h01;
ROM_MEM[4777] <= 8'h91;
ROM_MEM[4778] <= 8'h02;
ROM_MEM[4779] <= 8'h27;
ROM_MEM[4780] <= 8'h24;
ROM_MEM[4781] <= 8'h23;
ROM_MEM[4782] <= 8'h12;
ROM_MEM[4783] <= 8'h86;
ROM_MEM[4784] <= 8'h04;
ROM_MEM[4785] <= 8'h97;
ROM_MEM[4786] <= 8'hBD;
ROM_MEM[4787] <= 8'hA6;
ROM_MEM[4788] <= 8'h84;
ROM_MEM[4789] <= 8'h98;
ROM_MEM[4790] <= 8'h02;
ROM_MEM[4791] <= 8'hA7;
ROM_MEM[4792] <= 8'h84;
ROM_MEM[4793] <= 8'hBD;
ROM_MEM[4794] <= 8'h97;
ROM_MEM[4795] <= 8'hF2;
ROM_MEM[4796] <= 8'hBD;
ROM_MEM[4797] <= 8'hBD;
ROM_MEM[4798] <= 8'hFD;
ROM_MEM[4799] <= 8'h20;
ROM_MEM[4800] <= 8'h10;
ROM_MEM[4801] <= 8'h86;
ROM_MEM[4802] <= 8'h04;
ROM_MEM[4803] <= 8'h97;
ROM_MEM[4804] <= 8'hBD;
ROM_MEM[4805] <= 8'hA6;
ROM_MEM[4806] <= 8'h84;
ROM_MEM[4807] <= 8'h98;
ROM_MEM[4808] <= 8'h02;
ROM_MEM[4809] <= 8'hA7;
ROM_MEM[4810] <= 8'h84;
ROM_MEM[4811] <= 8'hBD;
ROM_MEM[4812] <= 8'h97;
ROM_MEM[4813] <= 8'hFC;
ROM_MEM[4814] <= 8'hBD;
ROM_MEM[4815] <= 8'hBD;
ROM_MEM[4816] <= 8'hFD;
ROM_MEM[4817] <= 8'h39;
ROM_MEM[4818] <= 8'h96;
ROM_MEM[4819] <= 8'hBC;
ROM_MEM[4820] <= 8'h27;
ROM_MEM[4821] <= 8'h0D;
ROM_MEM[4822] <= 8'hDC;
ROM_MEM[4823] <= 8'hCC;
ROM_MEM[4824] <= 8'h2B;
ROM_MEM[4825] <= 8'h07;
ROM_MEM[4826] <= 8'h86;
ROM_MEM[4827] <= 8'h04;
ROM_MEM[4828] <= 8'h97;
ROM_MEM[4829] <= 8'hBD;
ROM_MEM[4830] <= 8'hBD;
ROM_MEM[4831] <= 8'hAD;
ROM_MEM[4832] <= 8'h20;
ROM_MEM[4833] <= 8'h20;
ROM_MEM[4834] <= 8'h01;
ROM_MEM[4835] <= 8'h39;
ROM_MEM[4836] <= 8'hDC;
ROM_MEM[4837] <= 8'hC4;
ROM_MEM[4838] <= 8'h2B;
ROM_MEM[4839] <= 8'h10;
ROM_MEM[4840] <= 8'h10;
ROM_MEM[4841] <= 8'h93;
ROM_MEM[4842] <= 8'hC8;
ROM_MEM[4843] <= 8'h22;
ROM_MEM[4844] <= 8'h0B;
ROM_MEM[4845] <= 8'h93;
ROM_MEM[4846] <= 8'hD0;
ROM_MEM[4847] <= 8'h22;
ROM_MEM[4848] <= 8'h16;
ROM_MEM[4849] <= 8'h86;
ROM_MEM[4850] <= 8'h04;
ROM_MEM[4851] <= 8'h97;
ROM_MEM[4852] <= 8'hBD;
ROM_MEM[4853] <= 8'h7E;
ROM_MEM[4854] <= 8'h8A;
ROM_MEM[4855] <= 8'hCF;
ROM_MEM[4856] <= 8'hDC;
ROM_MEM[4857] <= 8'hC8;
ROM_MEM[4858] <= 8'h2B;
ROM_MEM[4859] <= 8'h0B;
ROM_MEM[4860] <= 8'h93;
ROM_MEM[4861] <= 8'hD0;
ROM_MEM[4862] <= 8'h22;
ROM_MEM[4863] <= 8'h07;
ROM_MEM[4864] <= 8'h86;
ROM_MEM[4865] <= 8'h04;
ROM_MEM[4866] <= 8'h97;
ROM_MEM[4867] <= 8'hBD;
ROM_MEM[4868] <= 8'h7E;
ROM_MEM[4869] <= 8'hA5;
ROM_MEM[4870] <= 8'h4B;
ROM_MEM[4871] <= 8'hDC;
ROM_MEM[4872] <= 8'hD0;
ROM_MEM[4873] <= 8'h2B;
ROM_MEM[4874] <= 8'h1F;
ROM_MEM[4875] <= 8'h86;
ROM_MEM[4876] <= 8'hFF;
ROM_MEM[4877] <= 8'h97;
ROM_MEM[4878] <= 8'hBD;
ROM_MEM[4879] <= 8'h86;
ROM_MEM[4880] <= 8'h0F;
ROM_MEM[4881] <= 8'hB7;
ROM_MEM[4882] <= 8'h4B;
ROM_MEM[4883] <= 8'h23;
ROM_MEM[4884] <= 8'h96;
ROM_MEM[4885] <= 8'hD0;
ROM_MEM[4886] <= 8'hC6;
ROM_MEM[4887] <= 8'h03;
ROM_MEM[4888] <= 8'h3D;
ROM_MEM[4889] <= 8'h10;
ROM_MEM[4890] <= 8'h83;
ROM_MEM[4891] <= 8'h00;
ROM_MEM[4892] <= 8'hE0;
ROM_MEM[4893] <= 8'h25;
ROM_MEM[4894] <= 8'h02;
ROM_MEM[4895] <= 8'hC6;
ROM_MEM[4896] <= 8'hE0;
ROM_MEM[4897] <= 8'hF7;
ROM_MEM[4898] <= 8'h4B;
ROM_MEM[4899] <= 8'h22;
ROM_MEM[4900] <= 8'hCC;
ROM_MEM[4901] <= 8'h66;
ROM_MEM[4902] <= 8'h80;
ROM_MEM[4903] <= 8'hFD;
ROM_MEM[4904] <= 8'h4B;
ROM_MEM[4905] <= 8'h20;
ROM_MEM[4906] <= 8'h39;
ROM_MEM[4907] <= 8'h96;
ROM_MEM[4908] <= 8'hBC;
ROM_MEM[4909] <= 8'h27;
ROM_MEM[4910] <= 8'h0E;
ROM_MEM[4911] <= 8'hDC;
ROM_MEM[4912] <= 8'hCC;
ROM_MEM[4913] <= 8'h2B;
ROM_MEM[4914] <= 8'h06;
ROM_MEM[4915] <= 8'h93;
ROM_MEM[4916] <= 8'hC4;
ROM_MEM[4917] <= 8'h25;
ROM_MEM[4918] <= 8'h07;
ROM_MEM[4919] <= 8'h20;
ROM_MEM[4920] <= 8'h0C;
ROM_MEM[4921] <= 8'h96;
ROM_MEM[4922] <= 8'hC4;
ROM_MEM[4923] <= 8'h2C;
ROM_MEM[4924] <= 8'h08;
ROM_MEM[4925] <= 8'h39;
ROM_MEM[4926] <= 8'h86;
ROM_MEM[4927] <= 8'h04;
ROM_MEM[4928] <= 8'h97;
ROM_MEM[4929] <= 8'hBD;
ROM_MEM[4930] <= 8'h7E;
ROM_MEM[4931] <= 8'hAD;
ROM_MEM[4932] <= 8'h20;
ROM_MEM[4933] <= 8'h86;
ROM_MEM[4934] <= 8'h04;
ROM_MEM[4935] <= 8'h97;
ROM_MEM[4936] <= 8'hBD;
ROM_MEM[4937] <= 8'h7E;
ROM_MEM[4938] <= 8'h8A;
ROM_MEM[4939] <= 8'hCF;
ROM_MEM[4940] <= 8'hB9;
ROM_MEM[4941] <= 8'h94;
ROM_MEM[4942] <= 8'hFF;
ROM_MEM[4943] <= 8'hFF;
ROM_MEM[4944] <= 8'hFF;
ROM_MEM[4945] <= 8'hFF;
ROM_MEM[4946] <= 8'hFF;
ROM_MEM[4947] <= 8'hFF;
ROM_MEM[4948] <= 8'hFF;
ROM_MEM[4949] <= 8'hFF;
ROM_MEM[4950] <= 8'hFF;
ROM_MEM[4951] <= 8'hFF;
ROM_MEM[4952] <= 8'hFF;
ROM_MEM[4953] <= 8'hFF;
ROM_MEM[4954] <= 8'hFF;
ROM_MEM[4955] <= 8'hFF;
ROM_MEM[4956] <= 8'hFF;
ROM_MEM[4957] <= 8'hFF;
ROM_MEM[4958] <= 8'hFF;
ROM_MEM[4959] <= 8'hFF;
ROM_MEM[4960] <= 8'hFF;
ROM_MEM[4961] <= 8'hFF;
ROM_MEM[4962] <= 8'hFF;
ROM_MEM[4963] <= 8'hFF;
ROM_MEM[4964] <= 8'hFF;
ROM_MEM[4965] <= 8'hFF;
ROM_MEM[4966] <= 8'hFF;
ROM_MEM[4967] <= 8'hFF;
ROM_MEM[4968] <= 8'hFF;
ROM_MEM[4969] <= 8'hFF;
ROM_MEM[4970] <= 8'hFF;
ROM_MEM[4971] <= 8'hFF;
ROM_MEM[4972] <= 8'hFF;
ROM_MEM[4973] <= 8'hFF;
ROM_MEM[4974] <= 8'hFF;
ROM_MEM[4975] <= 8'hFF;
ROM_MEM[4976] <= 8'hFF;
ROM_MEM[4977] <= 8'hFF;
ROM_MEM[4978] <= 8'hFF;
ROM_MEM[4979] <= 8'hFF;
ROM_MEM[4980] <= 8'hFF;
ROM_MEM[4981] <= 8'hFF;
ROM_MEM[4982] <= 8'hFF;
ROM_MEM[4983] <= 8'hFF;
ROM_MEM[4984] <= 8'hFF;
ROM_MEM[4985] <= 8'hFF;
ROM_MEM[4986] <= 8'hFF;
ROM_MEM[4987] <= 8'hFF;
ROM_MEM[4988] <= 8'hFF;
ROM_MEM[4989] <= 8'hFF;
ROM_MEM[4990] <= 8'hFF;
ROM_MEM[4991] <= 8'hFF;
ROM_MEM[4992] <= 8'hFF;
ROM_MEM[4993] <= 8'hFF;
ROM_MEM[4994] <= 8'hFF;
ROM_MEM[4995] <= 8'hFF;
ROM_MEM[4996] <= 8'hFF;
ROM_MEM[4997] <= 8'hFF;
ROM_MEM[4998] <= 8'hFF;
ROM_MEM[4999] <= 8'hFF;
ROM_MEM[5000] <= 8'hFF;
ROM_MEM[5001] <= 8'hFF;
ROM_MEM[5002] <= 8'hFF;
ROM_MEM[5003] <= 8'hFF;
ROM_MEM[5004] <= 8'hFF;
ROM_MEM[5005] <= 8'hFF;
ROM_MEM[5006] <= 8'hFF;
ROM_MEM[5007] <= 8'hFF;
ROM_MEM[5008] <= 8'hFF;
ROM_MEM[5009] <= 8'hFF;
ROM_MEM[5010] <= 8'hFF;
ROM_MEM[5011] <= 8'hFF;
ROM_MEM[5012] <= 8'hFF;
ROM_MEM[5013] <= 8'hFF;
ROM_MEM[5014] <= 8'hFF;
ROM_MEM[5015] <= 8'hFF;
ROM_MEM[5016] <= 8'hFF;
ROM_MEM[5017] <= 8'hFF;
ROM_MEM[5018] <= 8'hFF;
ROM_MEM[5019] <= 8'hFF;
ROM_MEM[5020] <= 8'hFF;
ROM_MEM[5021] <= 8'hFF;
ROM_MEM[5022] <= 8'hFF;
ROM_MEM[5023] <= 8'hFF;
ROM_MEM[5024] <= 8'hFF;
ROM_MEM[5025] <= 8'hFF;
ROM_MEM[5026] <= 8'hFF;
ROM_MEM[5027] <= 8'hFF;
ROM_MEM[5028] <= 8'hFF;
ROM_MEM[5029] <= 8'hFF;
ROM_MEM[5030] <= 8'hFF;
ROM_MEM[5031] <= 8'hFF;
ROM_MEM[5032] <= 8'hFF;
ROM_MEM[5033] <= 8'hFF;
ROM_MEM[5034] <= 8'hFF;
ROM_MEM[5035] <= 8'hFF;
ROM_MEM[5036] <= 8'hFF;
ROM_MEM[5037] <= 8'hFF;
ROM_MEM[5038] <= 8'hFF;
ROM_MEM[5039] <= 8'hFF;
ROM_MEM[5040] <= 8'hFF;
ROM_MEM[5041] <= 8'hFF;
ROM_MEM[5042] <= 8'h43;
ROM_MEM[5043] <= 8'h4F;
ROM_MEM[5044] <= 8'h50;
ROM_MEM[5045] <= 8'h59;
ROM_MEM[5046] <= 8'h52;
ROM_MEM[5047] <= 8'h49;
ROM_MEM[5048] <= 8'h47;
ROM_MEM[5049] <= 8'h48;
ROM_MEM[5050] <= 8'h54;
ROM_MEM[5051] <= 8'h20;
ROM_MEM[5052] <= 8'h31;
ROM_MEM[5053] <= 8'h39;
ROM_MEM[5054] <= 8'h38;
ROM_MEM[5055] <= 8'h33;
ROM_MEM[5056] <= 8'h20;
ROM_MEM[5057] <= 8'h41;
ROM_MEM[5058] <= 8'h54;
ROM_MEM[5059] <= 8'h41;
ROM_MEM[5060] <= 8'h52;
ROM_MEM[5061] <= 8'h49;
ROM_MEM[5062] <= 8'h04;
ROM_MEM[5063] <= 8'hBC;
ROM_MEM[5064] <= 8'h96;
ROM_MEM[5065] <= 8'hFA;
ROM_MEM[5066] <= 8'h5B;
ROM_MEM[5067] <= 8'h28;
ROM_MEM[5068] <= 8'h41;
ROM_MEM[5069] <= 8'h4C;
ROM_MEM[5070] <= 8'h4C;
ROM_MEM[5071] <= 8'h59;
ROM_MEM[5072] <= 8'h20;
ROM_MEM[5073] <= 8'h57;
ROM_MEM[5074] <= 8'h41;
ROM_MEM[5075] <= 8'h53;
ROM_MEM[5076] <= 8'h20;
ROM_MEM[5077] <= 8'h54;
ROM_MEM[5078] <= 8'h48;
ROM_MEM[5079] <= 8'h45;
ROM_MEM[5080] <= 8'h20;
ROM_MEM[5081] <= 8'h57;
ROM_MEM[5082] <= 8'h48;
ROM_MEM[5083] <= 8'h49;
ROM_MEM[5084] <= 8'h50;
ROM_MEM[5085] <= 8'h43;
ROM_MEM[5086] <= 8'h52;
ROM_MEM[5087] <= 8'h41;
ROM_MEM[5088] <= 8'h43;
ROM_MEM[5089] <= 8'h4B;
ROM_MEM[5090] <= 8'h45;
ROM_MEM[5091] <= 8'h52;
ROM_MEM[5092] <= 8'hB6;
ROM_MEM[5093] <= 8'h49;
ROM_MEM[5094] <= 8'hC0;
ROM_MEM[5095] <= 8'h81;
ROM_MEM[5096] <= 8'h03;
ROM_MEM[5097] <= 8'h25;
ROM_MEM[5098] <= 8'h05;
ROM_MEM[5099] <= 8'h86;
ROM_MEM[5100] <= 8'h00;
ROM_MEM[5101] <= 8'hB7;
ROM_MEM[5102] <= 8'h49;
ROM_MEM[5103] <= 8'hC0;
ROM_MEM[5104] <= 8'h86;
ROM_MEM[5105] <= 8'h01;
ROM_MEM[5106] <= 8'h97;
ROM_MEM[5107] <= 8'h9C;
ROM_MEM[5108] <= 8'h86;
ROM_MEM[5109] <= 8'h0B;
ROM_MEM[5110] <= 8'h97;
ROM_MEM[5111] <= 8'hDC;
ROM_MEM[5112] <= 8'h97;
ROM_MEM[5113] <= 8'h9D;
ROM_MEM[5114] <= 8'hBD;
ROM_MEM[5115] <= 8'hCD;
ROM_MEM[5116] <= 8'h38;
ROM_MEM[5117] <= 8'hBD;
ROM_MEM[5118] <= 8'hB4;
ROM_MEM[5119] <= 8'h3F;
ROM_MEM[5120] <= 8'h96;
ROM_MEM[5121] <= 8'h9D;
ROM_MEM[5122] <= 8'h97;
ROM_MEM[5123] <= 8'hDC;
ROM_MEM[5124] <= 8'hBD;
ROM_MEM[5125] <= 8'hCD;
ROM_MEM[5126] <= 8'h44;
ROM_MEM[5127] <= 8'hBD;
ROM_MEM[5128] <= 8'hB5;
ROM_MEM[5129] <= 8'h79;
ROM_MEM[5130] <= 8'h86;
ROM_MEM[5131] <= 8'h02;
ROM_MEM[5132] <= 8'h97;
ROM_MEM[5133] <= 8'h9C;
ROM_MEM[5134] <= 8'h86;
ROM_MEM[5135] <= 8'h0E;
ROM_MEM[5136] <= 8'h97;
ROM_MEM[5137] <= 8'hDC;
ROM_MEM[5138] <= 8'h97;
ROM_MEM[5139] <= 8'h9D;
ROM_MEM[5140] <= 8'hBD;
ROM_MEM[5141] <= 8'hCD;
ROM_MEM[5142] <= 8'h38;
ROM_MEM[5143] <= 8'hBD;
ROM_MEM[5144] <= 8'hB4;
ROM_MEM[5145] <= 8'h3F;
ROM_MEM[5146] <= 8'h96;
ROM_MEM[5147] <= 8'h9D;
ROM_MEM[5148] <= 8'h97;
ROM_MEM[5149] <= 8'hDC;
ROM_MEM[5150] <= 8'hBD;
ROM_MEM[5151] <= 8'hCD;
ROM_MEM[5152] <= 8'h44;
ROM_MEM[5153] <= 8'hBD;
ROM_MEM[5154] <= 8'hB5;
ROM_MEM[5155] <= 8'h79;
ROM_MEM[5156] <= 8'h86;
ROM_MEM[5157] <= 8'h03;
ROM_MEM[5158] <= 8'h97;
ROM_MEM[5159] <= 8'h9C;
ROM_MEM[5160] <= 8'h86;
ROM_MEM[5161] <= 8'h0C;
ROM_MEM[5162] <= 8'h97;
ROM_MEM[5163] <= 8'hDC;
ROM_MEM[5164] <= 8'h97;
ROM_MEM[5165] <= 8'h9D;
ROM_MEM[5166] <= 8'hBD;
ROM_MEM[5167] <= 8'hCD;
ROM_MEM[5168] <= 8'h38;
ROM_MEM[5169] <= 8'hBD;
ROM_MEM[5170] <= 8'hB4;
ROM_MEM[5171] <= 8'h3F;
ROM_MEM[5172] <= 8'h96;
ROM_MEM[5173] <= 8'h9D;
ROM_MEM[5174] <= 8'h97;
ROM_MEM[5175] <= 8'hDC;
ROM_MEM[5176] <= 8'hBD;
ROM_MEM[5177] <= 8'hCD;
ROM_MEM[5178] <= 8'h44;
ROM_MEM[5179] <= 8'hBD;
ROM_MEM[5180] <= 8'hB5;
ROM_MEM[5181] <= 8'h79;
ROM_MEM[5182] <= 8'h39;
ROM_MEM[5183] <= 8'h86;
ROM_MEM[5184] <= 8'h00;
ROM_MEM[5185] <= 8'hB7;
ROM_MEM[5186] <= 8'h49;
ROM_MEM[5187] <= 8'hBD;
ROM_MEM[5188] <= 8'hB6;
ROM_MEM[5189] <= 8'h49;
ROM_MEM[5190] <= 8'hC0;
ROM_MEM[5191] <= 8'hB7;
ROM_MEM[5192] <= 8'h49;
ROM_MEM[5193] <= 8'hBE;
ROM_MEM[5194] <= 8'h86;
ROM_MEM[5195] <= 8'h88;
ROM_MEM[5196] <= 8'hB7;
ROM_MEM[5197] <= 8'h49;
ROM_MEM[5198] <= 8'hC1;
ROM_MEM[5199] <= 8'hF6;
ROM_MEM[5200] <= 8'h50;
ROM_MEM[5201] <= 8'h40;
ROM_MEM[5202] <= 8'h54;
ROM_MEM[5203] <= 8'h54;
ROM_MEM[5204] <= 8'h54;
ROM_MEM[5205] <= 8'hC4;
ROM_MEM[5206] <= 8'h0F;
ROM_MEM[5207] <= 8'h8E;
ROM_MEM[5208] <= 8'h49;
ROM_MEM[5209] <= 8'h89;
ROM_MEM[5210] <= 8'h3A;
ROM_MEM[5211] <= 8'h9F;
ROM_MEM[5212] <= 8'h64;
ROM_MEM[5213] <= 8'hB6;
ROM_MEM[5214] <= 8'h50;
ROM_MEM[5215] <= 8'h40;
ROM_MEM[5216] <= 8'h84;
ROM_MEM[5217] <= 8'hF8;
ROM_MEM[5218] <= 8'h8B;
ROM_MEM[5219] <= 8'h04;
ROM_MEM[5220] <= 8'hC6;
ROM_MEM[5221] <= 8'h00;
ROM_MEM[5222] <= 8'hFD;
ROM_MEM[5223] <= 8'h50;
ROM_MEM[5224] <= 8'h78;
ROM_MEM[5225] <= 8'hCC;
ROM_MEM[5226] <= 8'hFC;
ROM_MEM[5227] <= 8'h00;
ROM_MEM[5228] <= 8'hFD;
ROM_MEM[5229] <= 8'h50;
ROM_MEM[5230] <= 8'h7A;
ROM_MEM[5231] <= 8'hCC;
ROM_MEM[5232] <= 8'hF2;
ROM_MEM[5233] <= 8'h00;
ROM_MEM[5234] <= 8'hFD;
ROM_MEM[5235] <= 8'h50;
ROM_MEM[5236] <= 8'h7C;
ROM_MEM[5237] <= 8'h9E;
ROM_MEM[5238] <= 8'h64;
ROM_MEM[5239] <= 8'h8C;
ROM_MEM[5240] <= 8'h49;
ROM_MEM[5241] <= 8'h99;
ROM_MEM[5242] <= 8'h25;
ROM_MEM[5243] <= 8'h03;
ROM_MEM[5244] <= 8'h30;
ROM_MEM[5245] <= 8'h88;
ROM_MEM[5246] <= 8'hF0;
ROM_MEM[5247] <= 8'hA6;
ROM_MEM[5248] <= 8'h80;
ROM_MEM[5249] <= 8'h9F;
ROM_MEM[5250] <= 8'h64;
ROM_MEM[5251] <= 8'h97;
ROM_MEM[5252] <= 8'h9E;
ROM_MEM[5253] <= 8'h84;
ROM_MEM[5254] <= 8'h03;
ROM_MEM[5255] <= 8'h91;
ROM_MEM[5256] <= 8'h9C;
ROM_MEM[5257] <= 8'h10;
ROM_MEM[5258] <= 8'h26;
ROM_MEM[5259] <= 8'h00;
ROM_MEM[5260] <= 8'h89;
ROM_MEM[5261] <= 8'h96;
ROM_MEM[5262] <= 8'h9D;
ROM_MEM[5263] <= 8'h97;
ROM_MEM[5264] <= 8'hDC;
ROM_MEM[5265] <= 8'hCC;
ROM_MEM[5266] <= 8'h00;
ROM_MEM[5267] <= 8'h0F;
ROM_MEM[5268] <= 8'hFD;
ROM_MEM[5269] <= 8'h47;
ROM_MEM[5270] <= 8'h01;
ROM_MEM[5271] <= 8'h86;
ROM_MEM[5272] <= 8'h67;
ROM_MEM[5273] <= 8'hBD;
ROM_MEM[5274] <= 8'hCD;
ROM_MEM[5275] <= 8'hBA;
ROM_MEM[5276] <= 8'h96;
ROM_MEM[5277] <= 8'h9C;
ROM_MEM[5278] <= 8'h81;
ROM_MEM[5279] <= 8'h02;
ROM_MEM[5280] <= 8'h26;
ROM_MEM[5281] <= 8'h13;
ROM_MEM[5282] <= 8'h7C;
ROM_MEM[5283] <= 8'h49;
ROM_MEM[5284] <= 8'hBD;
ROM_MEM[5285] <= 8'hF6;
ROM_MEM[5286] <= 8'h49;
ROM_MEM[5287] <= 8'hBE;
ROM_MEM[5288] <= 8'h58;
ROM_MEM[5289] <= 8'h8E;
ROM_MEM[5290] <= 8'hB6;
ROM_MEM[5291] <= 8'hB3;
ROM_MEM[5292] <= 8'hEC;
ROM_MEM[5293] <= 8'h85;
ROM_MEM[5294] <= 8'hED;
ROM_MEM[5295] <= 8'hA1;
ROM_MEM[5296] <= 8'hB6;
ROM_MEM[5297] <= 8'h49;
ROM_MEM[5298] <= 8'hC1;
ROM_MEM[5299] <= 8'hA7;
ROM_MEM[5300] <= 8'h3F;
ROM_MEM[5301] <= 8'hFC;
ROM_MEM[5302] <= 8'h50;
ROM_MEM[5303] <= 8'h78;
ROM_MEM[5304] <= 8'hB3;
ROM_MEM[5305] <= 8'h50;
ROM_MEM[5306] <= 8'h40;
ROM_MEM[5307] <= 8'h10;
ROM_MEM[5308] <= 8'h83;
ROM_MEM[5309] <= 8'h10;
ROM_MEM[5310] <= 8'h00;
ROM_MEM[5311] <= 8'h2E;
ROM_MEM[5312] <= 8'h4F;
ROM_MEM[5313] <= 8'h96;
ROM_MEM[5314] <= 8'h9D;
ROM_MEM[5315] <= 8'h81;
ROM_MEM[5316] <= 8'h0E;
ROM_MEM[5317] <= 8'h26;
ROM_MEM[5318] <= 8'h44;
ROM_MEM[5319] <= 8'hFC;
ROM_MEM[5320] <= 8'h50;
ROM_MEM[5321] <= 8'h00;
ROM_MEM[5322] <= 8'h83;
ROM_MEM[5323] <= 8'h00;
ROM_MEM[5324] <= 8'h00;
ROM_MEM[5325] <= 8'h2D;
ROM_MEM[5326] <= 8'h47;
ROM_MEM[5327] <= 8'hFC;
ROM_MEM[5328] <= 8'h50;
ROM_MEM[5329] <= 8'h42;
ROM_MEM[5330] <= 8'h2E;
ROM_MEM[5331] <= 8'h37;
ROM_MEM[5332] <= 8'hFC;
ROM_MEM[5333] <= 8'h50;
ROM_MEM[5334] <= 8'h7C;
ROM_MEM[5335] <= 8'hC3;
ROM_MEM[5336] <= 8'h02;
ROM_MEM[5337] <= 8'h00;
ROM_MEM[5338] <= 8'hB3;
ROM_MEM[5339] <= 8'h50;
ROM_MEM[5340] <= 8'h44;
ROM_MEM[5341] <= 8'h2D;
ROM_MEM[5342] <= 8'h2C;
ROM_MEM[5343] <= 8'h83;
ROM_MEM[5344] <= 8'h04;
ROM_MEM[5345] <= 8'h00;
ROM_MEM[5346] <= 8'h2E;
ROM_MEM[5347] <= 8'h27;
ROM_MEM[5348] <= 8'hFC;
ROM_MEM[5349] <= 8'h50;
ROM_MEM[5350] <= 8'h78;
ROM_MEM[5351] <= 8'hB3;
ROM_MEM[5352] <= 8'h50;
ROM_MEM[5353] <= 8'h40;
ROM_MEM[5354] <= 8'h83;
ROM_MEM[5355] <= 8'h04;
ROM_MEM[5356] <= 8'h00;
ROM_MEM[5357] <= 8'h22;
ROM_MEM[5358] <= 8'h1C;
ROM_MEM[5359] <= 8'h86;
ROM_MEM[5360] <= 8'h0F;
ROM_MEM[5361] <= 8'h97;
ROM_MEM[5362] <= 8'hDC;
ROM_MEM[5363] <= 8'h96;
ROM_MEM[5364] <= 8'h60;
ROM_MEM[5365] <= 8'h2D;
ROM_MEM[5366] <= 8'h06;
ROM_MEM[5367] <= 8'hBD;
ROM_MEM[5368] <= 8'h98;
ROM_MEM[5369] <= 8'h74;
ROM_MEM[5370] <= 8'hBD;
ROM_MEM[5371] <= 8'hBD;
ROM_MEM[5372] <= 8'hB2;
ROM_MEM[5373] <= 8'h96;
ROM_MEM[5374] <= 8'h63;
ROM_MEM[5375] <= 8'h26;
ROM_MEM[5376] <= 8'h0A;
ROM_MEM[5377] <= 8'h86;
ROM_MEM[5378] <= 8'h4E;
ROM_MEM[5379] <= 8'hF6;
ROM_MEM[5380] <= 8'h47;
ROM_MEM[5381] <= 8'h03;
ROM_MEM[5382] <= 8'h2A;
ROM_MEM[5383] <= 8'h01;
ROM_MEM[5384] <= 8'h40;
ROM_MEM[5385] <= 8'h97;
ROM_MEM[5386] <= 8'h63;
ROM_MEM[5387] <= 8'hBD;
ROM_MEM[5388] <= 8'hCD;
ROM_MEM[5389] <= 8'h5C;
ROM_MEM[5390] <= 8'h20;
ROM_MEM[5391] <= 8'h03;
ROM_MEM[5392] <= 8'hBD;
ROM_MEM[5393] <= 8'hCD;
ROM_MEM[5394] <= 8'h50;
ROM_MEM[5395] <= 8'hBD;
ROM_MEM[5396] <= 8'hCD;
ROM_MEM[5397] <= 8'h74;
ROM_MEM[5398] <= 8'hFC;
ROM_MEM[5399] <= 8'h50;
ROM_MEM[5400] <= 8'h7C;
ROM_MEM[5401] <= 8'hC3;
ROM_MEM[5402] <= 8'h04;
ROM_MEM[5403] <= 8'h00;
ROM_MEM[5404] <= 8'hFD;
ROM_MEM[5405] <= 8'h50;
ROM_MEM[5406] <= 8'h7C;
ROM_MEM[5407] <= 8'h96;
ROM_MEM[5408] <= 8'h9E;
ROM_MEM[5409] <= 8'h44;
ROM_MEM[5410] <= 8'h44;
ROM_MEM[5411] <= 8'h10;
ROM_MEM[5412] <= 8'h26;
ROM_MEM[5413] <= 8'hFF;
ROM_MEM[5414] <= 8'h5C;
ROM_MEM[5415] <= 8'h96;
ROM_MEM[5416] <= 8'h9C;
ROM_MEM[5417] <= 8'h81;
ROM_MEM[5418] <= 8'h02;
ROM_MEM[5419] <= 8'h26;
ROM_MEM[5420] <= 8'h38;
ROM_MEM[5421] <= 8'h9E;
ROM_MEM[5422] <= 8'h64;
ROM_MEM[5423] <= 8'hA6;
ROM_MEM[5424] <= 8'h89;
ROM_MEM[5425] <= 8'h00;
ROM_MEM[5426] <= 8'h0F;
ROM_MEM[5427] <= 8'h48;
ROM_MEM[5428] <= 8'h24;
ROM_MEM[5429] <= 8'h07;
ROM_MEM[5430] <= 8'h2B;
ROM_MEM[5431] <= 8'h05;
ROM_MEM[5432] <= 8'h7C;
ROM_MEM[5433] <= 8'h49;
ROM_MEM[5434] <= 8'hBD;
ROM_MEM[5435] <= 8'h20;
ROM_MEM[5436] <= 8'h03;
ROM_MEM[5437] <= 8'h48;
ROM_MEM[5438] <= 8'h26;
ROM_MEM[5439] <= 8'hF3;
ROM_MEM[5440] <= 8'hB6;
ROM_MEM[5441] <= 8'h49;
ROM_MEM[5442] <= 8'hBD;
ROM_MEM[5443] <= 8'h27;
ROM_MEM[5444] <= 8'h20;
ROM_MEM[5445] <= 8'hB6;
ROM_MEM[5446] <= 8'h49;
ROM_MEM[5447] <= 8'hBE;
ROM_MEM[5448] <= 8'h4C;
ROM_MEM[5449] <= 8'h81;
ROM_MEM[5450] <= 8'h03;
ROM_MEM[5451] <= 8'h25;
ROM_MEM[5452] <= 8'h02;
ROM_MEM[5453] <= 8'h86;
ROM_MEM[5454] <= 8'h00;
ROM_MEM[5455] <= 8'hB7;
ROM_MEM[5456] <= 8'h49;
ROM_MEM[5457] <= 8'hBE;
ROM_MEM[5458] <= 8'hB6;
ROM_MEM[5459] <= 8'h49;
ROM_MEM[5460] <= 8'hC1;
ROM_MEM[5461] <= 8'h80;
ROM_MEM[5462] <= 8'h08;
ROM_MEM[5463] <= 8'h81;
ROM_MEM[5464] <= 8'h40;
ROM_MEM[5465] <= 8'h24;
ROM_MEM[5466] <= 8'h02;
ROM_MEM[5467] <= 8'h86;
ROM_MEM[5468] <= 8'h40;
ROM_MEM[5469] <= 8'hB7;
ROM_MEM[5470] <= 8'h49;
ROM_MEM[5471] <= 8'hC1;
ROM_MEM[5472] <= 8'h86;
ROM_MEM[5473] <= 8'h00;
ROM_MEM[5474] <= 8'hB7;
ROM_MEM[5475] <= 8'h49;
ROM_MEM[5476] <= 8'hBD;
ROM_MEM[5477] <= 8'hFC;
ROM_MEM[5478] <= 8'h50;
ROM_MEM[5479] <= 8'h78;
ROM_MEM[5480] <= 8'hC3;
ROM_MEM[5481] <= 8'h08;
ROM_MEM[5482] <= 8'h00;
ROM_MEM[5483] <= 8'hFD;
ROM_MEM[5484] <= 8'h50;
ROM_MEM[5485] <= 8'h78;
ROM_MEM[5486] <= 8'hB3;
ROM_MEM[5487] <= 8'h50;
ROM_MEM[5488] <= 8'h40;
ROM_MEM[5489] <= 8'h83;
ROM_MEM[5490] <= 8'h70;
ROM_MEM[5491] <= 8'h00;
ROM_MEM[5492] <= 8'h10;
ROM_MEM[5493] <= 8'h25;
ROM_MEM[5494] <= 8'hFE;
ROM_MEM[5495] <= 8'hF7;
ROM_MEM[5496] <= 8'h39;
ROM_MEM[5497] <= 8'h86;
ROM_MEM[5498] <= 8'h00;
ROM_MEM[5499] <= 8'hB7;
ROM_MEM[5500] <= 8'h49;
ROM_MEM[5501] <= 8'hBD;
ROM_MEM[5502] <= 8'hB6;
ROM_MEM[5503] <= 8'h49;
ROM_MEM[5504] <= 8'hC0;
ROM_MEM[5505] <= 8'hB7;
ROM_MEM[5506] <= 8'h49;
ROM_MEM[5507] <= 8'hBE;
ROM_MEM[5508] <= 8'h86;
ROM_MEM[5509] <= 8'h88;
ROM_MEM[5510] <= 8'hB7;
ROM_MEM[5511] <= 8'h49;
ROM_MEM[5512] <= 8'hC1;
ROM_MEM[5513] <= 8'hF6;
ROM_MEM[5514] <= 8'h50;
ROM_MEM[5515] <= 8'h40;
ROM_MEM[5516] <= 8'h54;
ROM_MEM[5517] <= 8'h54;
ROM_MEM[5518] <= 8'h54;
ROM_MEM[5519] <= 8'hC4;
ROM_MEM[5520] <= 8'h0F;
ROM_MEM[5521] <= 8'h8E;
ROM_MEM[5522] <= 8'h49;
ROM_MEM[5523] <= 8'h99;
ROM_MEM[5524] <= 8'h3A;
ROM_MEM[5525] <= 8'h9F;
ROM_MEM[5526] <= 8'h64;
ROM_MEM[5527] <= 8'hB6;
ROM_MEM[5528] <= 8'h50;
ROM_MEM[5529] <= 8'h40;
ROM_MEM[5530] <= 8'h84;
ROM_MEM[5531] <= 8'hF8;
ROM_MEM[5532] <= 8'h8B;
ROM_MEM[5533] <= 8'h04;
ROM_MEM[5534] <= 8'hC6;
ROM_MEM[5535] <= 8'h00;
ROM_MEM[5536] <= 8'hFD;
ROM_MEM[5537] <= 8'h50;
ROM_MEM[5538] <= 8'h78;
ROM_MEM[5539] <= 8'hCC;
ROM_MEM[5540] <= 8'h04;
ROM_MEM[5541] <= 8'h00;
ROM_MEM[5542] <= 8'hFD;
ROM_MEM[5543] <= 8'h50;
ROM_MEM[5544] <= 8'h7A;
ROM_MEM[5545] <= 8'hCC;
ROM_MEM[5546] <= 8'hF2;
ROM_MEM[5547] <= 8'h00;
ROM_MEM[5548] <= 8'hFD;
ROM_MEM[5549] <= 8'h50;
ROM_MEM[5550] <= 8'h7C;
ROM_MEM[5551] <= 8'h9E;
ROM_MEM[5552] <= 8'h64;
ROM_MEM[5553] <= 8'h8C;
ROM_MEM[5554] <= 8'h49;
ROM_MEM[5555] <= 8'hA9;
ROM_MEM[5556] <= 8'h25;
ROM_MEM[5557] <= 8'h03;
ROM_MEM[5558] <= 8'h30;
ROM_MEM[5559] <= 8'h88;
ROM_MEM[5560] <= 8'hF0;
ROM_MEM[5561] <= 8'hA6;
ROM_MEM[5562] <= 8'h80;
ROM_MEM[5563] <= 8'h9F;
ROM_MEM[5564] <= 8'h64;
ROM_MEM[5565] <= 8'h97;
ROM_MEM[5566] <= 8'h9E;
ROM_MEM[5567] <= 8'h84;
ROM_MEM[5568] <= 8'h03;
ROM_MEM[5569] <= 8'h91;
ROM_MEM[5570] <= 8'h9C;
ROM_MEM[5571] <= 8'h10;
ROM_MEM[5572] <= 8'h26;
ROM_MEM[5573] <= 8'h00;
ROM_MEM[5574] <= 8'h89;
ROM_MEM[5575] <= 8'h96;
ROM_MEM[5576] <= 8'h9D;
ROM_MEM[5577] <= 8'h97;
ROM_MEM[5578] <= 8'hDC;
ROM_MEM[5579] <= 8'hCC;
ROM_MEM[5580] <= 8'h00;
ROM_MEM[5581] <= 8'h0F;
ROM_MEM[5582] <= 8'hFD;
ROM_MEM[5583] <= 8'h47;
ROM_MEM[5584] <= 8'h01;
ROM_MEM[5585] <= 8'h86;
ROM_MEM[5586] <= 8'h67;
ROM_MEM[5587] <= 8'hBD;
ROM_MEM[5588] <= 8'hCD;
ROM_MEM[5589] <= 8'hBA;
ROM_MEM[5590] <= 8'h96;
ROM_MEM[5591] <= 8'h9C;
ROM_MEM[5592] <= 8'h81;
ROM_MEM[5593] <= 8'h02;
ROM_MEM[5594] <= 8'h26;
ROM_MEM[5595] <= 8'h13;
ROM_MEM[5596] <= 8'h7C;
ROM_MEM[5597] <= 8'h49;
ROM_MEM[5598] <= 8'hBD;
ROM_MEM[5599] <= 8'hF6;
ROM_MEM[5600] <= 8'h49;
ROM_MEM[5601] <= 8'hBE;
ROM_MEM[5602] <= 8'h58;
ROM_MEM[5603] <= 8'h8E;
ROM_MEM[5604] <= 8'hB6;
ROM_MEM[5605] <= 8'hB3;
ROM_MEM[5606] <= 8'hEC;
ROM_MEM[5607] <= 8'h85;
ROM_MEM[5608] <= 8'hED;
ROM_MEM[5609] <= 8'hA1;
ROM_MEM[5610] <= 8'hB6;
ROM_MEM[5611] <= 8'h49;
ROM_MEM[5612] <= 8'hC1;
ROM_MEM[5613] <= 8'hA7;
ROM_MEM[5614] <= 8'h3F;
ROM_MEM[5615] <= 8'hFC;
ROM_MEM[5616] <= 8'h50;
ROM_MEM[5617] <= 8'h78;
ROM_MEM[5618] <= 8'hB3;
ROM_MEM[5619] <= 8'h50;
ROM_MEM[5620] <= 8'h40;
ROM_MEM[5621] <= 8'h10;
ROM_MEM[5622] <= 8'h83;
ROM_MEM[5623] <= 8'h10;
ROM_MEM[5624] <= 8'h00;
ROM_MEM[5625] <= 8'h2E;
ROM_MEM[5626] <= 8'h4F;
ROM_MEM[5627] <= 8'h96;
ROM_MEM[5628] <= 8'h9D;
ROM_MEM[5629] <= 8'h81;
ROM_MEM[5630] <= 8'h0E;
ROM_MEM[5631] <= 8'h26;
ROM_MEM[5632] <= 8'h44;
ROM_MEM[5633] <= 8'hFC;
ROM_MEM[5634] <= 8'h50;
ROM_MEM[5635] <= 8'h00;
ROM_MEM[5636] <= 8'h83;
ROM_MEM[5637] <= 8'h00;
ROM_MEM[5638] <= 8'h00;
ROM_MEM[5639] <= 8'h2D;
ROM_MEM[5640] <= 8'h47;
ROM_MEM[5641] <= 8'hFC;
ROM_MEM[5642] <= 8'h50;
ROM_MEM[5643] <= 8'h42;
ROM_MEM[5644] <= 8'h2D;
ROM_MEM[5645] <= 8'h37;
ROM_MEM[5646] <= 8'hFC;
ROM_MEM[5647] <= 8'h50;
ROM_MEM[5648] <= 8'h7C;
ROM_MEM[5649] <= 8'hC3;
ROM_MEM[5650] <= 8'h02;
ROM_MEM[5651] <= 8'h00;
ROM_MEM[5652] <= 8'hB3;
ROM_MEM[5653] <= 8'h50;
ROM_MEM[5654] <= 8'h44;
ROM_MEM[5655] <= 8'h2D;
ROM_MEM[5656] <= 8'h2C;
ROM_MEM[5657] <= 8'h83;
ROM_MEM[5658] <= 8'h04;
ROM_MEM[5659] <= 8'h00;
ROM_MEM[5660] <= 8'h2E;
ROM_MEM[5661] <= 8'h27;
ROM_MEM[5662] <= 8'hFC;
ROM_MEM[5663] <= 8'h50;
ROM_MEM[5664] <= 8'h78;
ROM_MEM[5665] <= 8'hB3;
ROM_MEM[5666] <= 8'h50;
ROM_MEM[5667] <= 8'h40;
ROM_MEM[5668] <= 8'h83;
ROM_MEM[5669] <= 8'h04;
ROM_MEM[5670] <= 8'h00;
ROM_MEM[5671] <= 8'h22;
ROM_MEM[5672] <= 8'h1C;
ROM_MEM[5673] <= 8'h86;
ROM_MEM[5674] <= 8'h0F;
ROM_MEM[5675] <= 8'h97;
ROM_MEM[5676] <= 8'hDC;
ROM_MEM[5677] <= 8'h96;
ROM_MEM[5678] <= 8'h60;
ROM_MEM[5679] <= 8'h2D;
ROM_MEM[5680] <= 8'h06;
ROM_MEM[5681] <= 8'hBD;
ROM_MEM[5682] <= 8'h98;
ROM_MEM[5683] <= 8'h74;
ROM_MEM[5684] <= 8'hBD;
ROM_MEM[5685] <= 8'hBD;
ROM_MEM[5686] <= 8'hB2;
ROM_MEM[5687] <= 8'h96;
ROM_MEM[5688] <= 8'h63;
ROM_MEM[5689] <= 8'h26;
ROM_MEM[5690] <= 8'h0A;
ROM_MEM[5691] <= 8'h86;
ROM_MEM[5692] <= 8'h4E;
ROM_MEM[5693] <= 8'hF6;
ROM_MEM[5694] <= 8'h47;
ROM_MEM[5695] <= 8'h03;
ROM_MEM[5696] <= 8'h2A;
ROM_MEM[5697] <= 8'h01;
ROM_MEM[5698] <= 8'h40;
ROM_MEM[5699] <= 8'h97;
ROM_MEM[5700] <= 8'h63;
ROM_MEM[5701] <= 8'hBD;
ROM_MEM[5702] <= 8'hCD;
ROM_MEM[5703] <= 8'h5C;
ROM_MEM[5704] <= 8'h20;
ROM_MEM[5705] <= 8'h03;
ROM_MEM[5706] <= 8'hBD;
ROM_MEM[5707] <= 8'hCD;
ROM_MEM[5708] <= 8'h50;
ROM_MEM[5709] <= 8'hBD;
ROM_MEM[5710] <= 8'hCD;
ROM_MEM[5711] <= 8'h74;
ROM_MEM[5712] <= 8'hFC;
ROM_MEM[5713] <= 8'h50;
ROM_MEM[5714] <= 8'h7C;
ROM_MEM[5715] <= 8'hC3;
ROM_MEM[5716] <= 8'h04;
ROM_MEM[5717] <= 8'h00;
ROM_MEM[5718] <= 8'hFD;
ROM_MEM[5719] <= 8'h50;
ROM_MEM[5720] <= 8'h7C;
ROM_MEM[5721] <= 8'h96;
ROM_MEM[5722] <= 8'h9E;
ROM_MEM[5723] <= 8'h44;
ROM_MEM[5724] <= 8'h44;
ROM_MEM[5725] <= 8'h10;
ROM_MEM[5726] <= 8'h26;
ROM_MEM[5727] <= 8'hFF;
ROM_MEM[5728] <= 8'h5C;
ROM_MEM[5729] <= 8'h96;
ROM_MEM[5730] <= 8'h9C;
ROM_MEM[5731] <= 8'h81;
ROM_MEM[5732] <= 8'h02;
ROM_MEM[5733] <= 8'h26;
ROM_MEM[5734] <= 8'h38;
ROM_MEM[5735] <= 8'h9E;
ROM_MEM[5736] <= 8'h64;
ROM_MEM[5737] <= 8'hA6;
ROM_MEM[5738] <= 8'h89;
ROM_MEM[5739] <= 8'hFF;
ROM_MEM[5740] <= 8'hEF;
ROM_MEM[5741] <= 8'h48;
ROM_MEM[5742] <= 8'h24;
ROM_MEM[5743] <= 8'h07;
ROM_MEM[5744] <= 8'h2B;
ROM_MEM[5745] <= 8'h05;
ROM_MEM[5746] <= 8'h7C;
ROM_MEM[5747] <= 8'h49;
ROM_MEM[5748] <= 8'hBD;
ROM_MEM[5749] <= 8'h20;
ROM_MEM[5750] <= 8'h03;
ROM_MEM[5751] <= 8'h48;
ROM_MEM[5752] <= 8'h26;
ROM_MEM[5753] <= 8'hF3;
ROM_MEM[5754] <= 8'hB6;
ROM_MEM[5755] <= 8'h49;
ROM_MEM[5756] <= 8'hBD;
ROM_MEM[5757] <= 8'h27;
ROM_MEM[5758] <= 8'h20;
ROM_MEM[5759] <= 8'hB6;
ROM_MEM[5760] <= 8'h49;
ROM_MEM[5761] <= 8'hBE;
ROM_MEM[5762] <= 8'h4C;
ROM_MEM[5763] <= 8'h81;
ROM_MEM[5764] <= 8'h03;
ROM_MEM[5765] <= 8'h25;
ROM_MEM[5766] <= 8'h02;
ROM_MEM[5767] <= 8'h86;
ROM_MEM[5768] <= 8'h00;
ROM_MEM[5769] <= 8'hB7;
ROM_MEM[5770] <= 8'h49;
ROM_MEM[5771] <= 8'hBE;
ROM_MEM[5772] <= 8'hB6;
ROM_MEM[5773] <= 8'h49;
ROM_MEM[5774] <= 8'hC1;
ROM_MEM[5775] <= 8'h80;
ROM_MEM[5776] <= 8'h08;
ROM_MEM[5777] <= 8'h81;
ROM_MEM[5778] <= 8'h40;
ROM_MEM[5779] <= 8'h24;
ROM_MEM[5780] <= 8'h02;
ROM_MEM[5781] <= 8'h86;
ROM_MEM[5782] <= 8'h40;
ROM_MEM[5783] <= 8'hB7;
ROM_MEM[5784] <= 8'h49;
ROM_MEM[5785] <= 8'hC1;
ROM_MEM[5786] <= 8'h86;
ROM_MEM[5787] <= 8'h00;
ROM_MEM[5788] <= 8'hB7;
ROM_MEM[5789] <= 8'h49;
ROM_MEM[5790] <= 8'hBD;
ROM_MEM[5791] <= 8'hFC;
ROM_MEM[5792] <= 8'h50;
ROM_MEM[5793] <= 8'h78;
ROM_MEM[5794] <= 8'hC3;
ROM_MEM[5795] <= 8'h08;
ROM_MEM[5796] <= 8'h00;
ROM_MEM[5797] <= 8'hFD;
ROM_MEM[5798] <= 8'h50;
ROM_MEM[5799] <= 8'h78;
ROM_MEM[5800] <= 8'hB3;
ROM_MEM[5801] <= 8'h50;
ROM_MEM[5802] <= 8'h40;
ROM_MEM[5803] <= 8'h83;
ROM_MEM[5804] <= 8'h70;
ROM_MEM[5805] <= 8'h00;
ROM_MEM[5806] <= 8'h10;
ROM_MEM[5807] <= 8'h25;
ROM_MEM[5808] <= 8'hFE;
ROM_MEM[5809] <= 8'hF7;
ROM_MEM[5810] <= 8'h39;
ROM_MEM[5811] <= 8'h66;
ROM_MEM[5812] <= 8'h80;
ROM_MEM[5813] <= 8'h63;
ROM_MEM[5814] <= 8'h80;
ROM_MEM[5815] <= 8'h65;
ROM_MEM[5816] <= 8'h80;
ROM_MEM[5817] <= 8'hBD;
ROM_MEM[5818] <= 8'hB6;
ROM_MEM[5819] <= 8'hC7;
ROM_MEM[5820] <= 8'hBD;
ROM_MEM[5821] <= 8'hB6;
ROM_MEM[5822] <= 8'hD7;
ROM_MEM[5823] <= 8'h39;
ROM_MEM[5824] <= 8'hBD;
ROM_MEM[5825] <= 8'hB6;
ROM_MEM[5826] <= 8'hCC;
ROM_MEM[5827] <= 8'hBD;
ROM_MEM[5828] <= 8'hB6;
ROM_MEM[5829] <= 8'hD7;
ROM_MEM[5830] <= 8'h39;
ROM_MEM[5831] <= 8'hCC;
ROM_MEM[5832] <= 8'h63;
ROM_MEM[5833] <= 8'h80;
ROM_MEM[5834] <= 8'hED;
ROM_MEM[5835] <= 8'hA1;
ROM_MEM[5836] <= 8'hCC;
ROM_MEM[5837] <= 8'hA0;
ROM_MEM[5838] <= 8'h12;
ROM_MEM[5839] <= 8'hED;
ROM_MEM[5840] <= 8'hA1;
ROM_MEM[5841] <= 8'hFC;
ROM_MEM[5842] <= 8'h32;
ROM_MEM[5843] <= 8'hFE;
ROM_MEM[5844] <= 8'hED;
ROM_MEM[5845] <= 8'hA1;
ROM_MEM[5846] <= 8'h39;
ROM_MEM[5847] <= 8'h96;
ROM_MEM[5848] <= 8'h7D;
ROM_MEM[5849] <= 8'h2A;
ROM_MEM[5850] <= 8'h01;
ROM_MEM[5851] <= 8'h40;
ROM_MEM[5852] <= 8'hC6;
ROM_MEM[5853] <= 8'h6E;
ROM_MEM[5854] <= 8'h3D;
ROM_MEM[5855] <= 8'hD6;
ROM_MEM[5856] <= 8'h7D;
ROM_MEM[5857] <= 8'h2A;
ROM_MEM[5858] <= 8'h01;
ROM_MEM[5859] <= 8'h40;
ROM_MEM[5860] <= 8'h1F;
ROM_MEM[5861] <= 8'h89;
ROM_MEM[5862] <= 8'h1D;
ROM_MEM[5863] <= 8'hFD;
ROM_MEM[5864] <= 8'h4B;
ROM_MEM[5865] <= 8'h1C;
ROM_MEM[5866] <= 8'h84;
ROM_MEM[5867] <= 8'h1F;
ROM_MEM[5868] <= 8'hED;
ROM_MEM[5869] <= 8'h22;
ROM_MEM[5870] <= 8'hED;
ROM_MEM[5871] <= 8'h28;
ROM_MEM[5872] <= 8'hED;
ROM_MEM[5873] <= 8'h2E;
ROM_MEM[5874] <= 8'hED;
ROM_MEM[5875] <= 8'hA8;
ROM_MEM[5876] <= 8'h14;
ROM_MEM[5877] <= 8'hED;
ROM_MEM[5878] <= 8'hA8;
ROM_MEM[5879] <= 8'h1A;
ROM_MEM[5880] <= 8'h96;
ROM_MEM[5881] <= 8'h7F;
ROM_MEM[5882] <= 8'h2A;
ROM_MEM[5883] <= 8'h01;
ROM_MEM[5884] <= 8'h40;
ROM_MEM[5885] <= 8'hC6;
ROM_MEM[5886] <= 8'h50;
ROM_MEM[5887] <= 8'h3D;
ROM_MEM[5888] <= 8'hD6;
ROM_MEM[5889] <= 8'h7F;
ROM_MEM[5890] <= 8'h2A;
ROM_MEM[5891] <= 8'h01;
ROM_MEM[5892] <= 8'h40;
ROM_MEM[5893] <= 8'h1F;
ROM_MEM[5894] <= 8'h89;
ROM_MEM[5895] <= 8'h1D;
ROM_MEM[5896] <= 8'hFD;
ROM_MEM[5897] <= 8'h4B;
ROM_MEM[5898] <= 8'h1E;
ROM_MEM[5899] <= 8'h84;
ROM_MEM[5900] <= 8'h1F;
ROM_MEM[5901] <= 8'hED;
ROM_MEM[5902] <= 8'hA4;
ROM_MEM[5903] <= 8'hED;
ROM_MEM[5904] <= 8'h26;
ROM_MEM[5905] <= 8'hED;
ROM_MEM[5906] <= 8'h2C;
ROM_MEM[5907] <= 8'hED;
ROM_MEM[5908] <= 8'hA8;
ROM_MEM[5909] <= 8'h12;
ROM_MEM[5910] <= 8'hED;
ROM_MEM[5911] <= 8'hA8;
ROM_MEM[5912] <= 8'h18;
ROM_MEM[5913] <= 8'hCC;
ROM_MEM[5914] <= 8'hBA;
ROM_MEM[5915] <= 8'hAC;
ROM_MEM[5916] <= 8'hED;
ROM_MEM[5917] <= 8'h24;
ROM_MEM[5918] <= 8'hCC;
ROM_MEM[5919] <= 8'hBA;
ROM_MEM[5920] <= 8'h0D;
ROM_MEM[5921] <= 8'hED;
ROM_MEM[5922] <= 8'h2A;
ROM_MEM[5923] <= 8'hCC;
ROM_MEM[5924] <= 8'hBB;
ROM_MEM[5925] <= 8'h33;
ROM_MEM[5926] <= 8'hED;
ROM_MEM[5927] <= 8'hA8;
ROM_MEM[5928] <= 8'h10;
ROM_MEM[5929] <= 8'hCC;
ROM_MEM[5930] <= 8'hBA;
ROM_MEM[5931] <= 8'hE6;
ROM_MEM[5932] <= 8'hED;
ROM_MEM[5933] <= 8'hA8;
ROM_MEM[5934] <= 8'h16;
ROM_MEM[5935] <= 8'hCC;
ROM_MEM[5936] <= 8'hBA;
ROM_MEM[5937] <= 8'h5A;
ROM_MEM[5938] <= 8'hED;
ROM_MEM[5939] <= 8'hA8;
ROM_MEM[5940] <= 8'h1C;
ROM_MEM[5941] <= 8'h31;
ROM_MEM[5942] <= 8'hA8;
ROM_MEM[5943] <= 8'h1E;
ROM_MEM[5944] <= 8'h39;
ROM_MEM[5945] <= 8'h86;
ROM_MEM[5946] <= 8'h00;
ROM_MEM[5947] <= 8'hA7;
ROM_MEM[5948] <= 8'h03;
ROM_MEM[5949] <= 8'hBD;
ROM_MEM[5950] <= 8'h8E;
ROM_MEM[5951] <= 8'h1C;
ROM_MEM[5952] <= 8'h34;
ROM_MEM[5953] <= 8'h50;
ROM_MEM[5954] <= 8'hBD;
ROM_MEM[5955] <= 8'hB7;
ROM_MEM[5956] <= 8'h6C;
ROM_MEM[5957] <= 8'h35;
ROM_MEM[5958] <= 8'h50;
ROM_MEM[5959] <= 8'h39;
ROM_MEM[5960] <= 8'hB9;
ROM_MEM[5961] <= 8'hC0;
ROM_MEM[5962] <= 8'hB9;
ROM_MEM[5963] <= 8'hC0;
ROM_MEM[5964] <= 8'hB9;
ROM_MEM[5965] <= 8'hC0;
ROM_MEM[5966] <= 8'hB9;
ROM_MEM[5967] <= 8'hC0;
ROM_MEM[5968] <= 8'hB9;
ROM_MEM[5969] <= 8'hC0;
ROM_MEM[5970] <= 8'hB9;
ROM_MEM[5971] <= 8'hC0;
ROM_MEM[5972] <= 8'hB9;
ROM_MEM[5973] <= 8'hF9;
ROM_MEM[5974] <= 8'hB9;
ROM_MEM[5975] <= 8'hF9;
ROM_MEM[5976] <= 8'hB9;
ROM_MEM[5977] <= 8'hF9;
ROM_MEM[5978] <= 8'hBA;
ROM_MEM[5979] <= 8'hA0;
ROM_MEM[5980] <= 8'hBA;
ROM_MEM[5981] <= 8'hA4;
ROM_MEM[5982] <= 8'hBA;
ROM_MEM[5983] <= 8'hA8;
ROM_MEM[5984] <= 8'hBA;
ROM_MEM[5985] <= 8'hAC;
ROM_MEM[5986] <= 8'hBA;
ROM_MEM[5987] <= 8'hB0;
ROM_MEM[5988] <= 8'hBA;
ROM_MEM[5989] <= 8'hB4;
ROM_MEM[5990] <= 8'hBB;
ROM_MEM[5991] <= 8'h1A;
ROM_MEM[5992] <= 8'hBB;
ROM_MEM[5993] <= 8'h1E;
ROM_MEM[5994] <= 8'hBB;
ROM_MEM[5995] <= 8'h16;
ROM_MEM[5996] <= 8'hEE;
ROM_MEM[5997] <= 8'h84;
ROM_MEM[5998] <= 8'hBD;
ROM_MEM[5999] <= 8'hB9;
ROM_MEM[6000] <= 8'h48;
ROM_MEM[6001] <= 8'h86;
ROM_MEM[6002] <= 8'h06;
ROM_MEM[6003] <= 8'hA7;
ROM_MEM[6004] <= 8'h0C;
ROM_MEM[6005] <= 8'h86;
ROM_MEM[6006] <= 8'h18;
ROM_MEM[6007] <= 8'hA7;
ROM_MEM[6008] <= 8'h0D;
ROM_MEM[6009] <= 8'hCC;
ROM_MEM[6010] <= 8'h00;
ROM_MEM[6011] <= 8'h00;
ROM_MEM[6012] <= 8'hA3;
ROM_MEM[6013] <= 8'h52;
ROM_MEM[6014] <= 8'hBD;
ROM_MEM[6015] <= 8'hCD;
ROM_MEM[6016] <= 8'h9C;
ROM_MEM[6017] <= 8'hED;
ROM_MEM[6018] <= 8'h06;
ROM_MEM[6019] <= 8'hE3;
ROM_MEM[6020] <= 8'h48;
ROM_MEM[6021] <= 8'hED;
ROM_MEM[6022] <= 8'h84;
ROM_MEM[6023] <= 8'hCC;
ROM_MEM[6024] <= 8'h00;
ROM_MEM[6025] <= 8'h00;
ROM_MEM[6026] <= 8'hA3;
ROM_MEM[6027] <= 8'h5A;
ROM_MEM[6028] <= 8'hBD;
ROM_MEM[6029] <= 8'hCD;
ROM_MEM[6030] <= 8'h9C;
ROM_MEM[6031] <= 8'hED;
ROM_MEM[6032] <= 8'h08;
ROM_MEM[6033] <= 8'hE3;
ROM_MEM[6034] <= 8'h4A;
ROM_MEM[6035] <= 8'hED;
ROM_MEM[6036] <= 8'h02;
ROM_MEM[6037] <= 8'hCC;
ROM_MEM[6038] <= 8'h00;
ROM_MEM[6039] <= 8'h00;
ROM_MEM[6040] <= 8'hA3;
ROM_MEM[6041] <= 8'h42;
ROM_MEM[6042] <= 8'hBD;
ROM_MEM[6043] <= 8'hCD;
ROM_MEM[6044] <= 8'h9C;
ROM_MEM[6045] <= 8'hED;
ROM_MEM[6046] <= 8'h0A;
ROM_MEM[6047] <= 8'hE3;
ROM_MEM[6048] <= 8'h4C;
ROM_MEM[6049] <= 8'hED;
ROM_MEM[6050] <= 8'h04;
ROM_MEM[6051] <= 8'hBD;
ROM_MEM[6052] <= 8'hB8;
ROM_MEM[6053] <= 8'h3F;
ROM_MEM[6054] <= 8'hBD;
ROM_MEM[6055] <= 8'hB9;
ROM_MEM[6056] <= 8'h48;
ROM_MEM[6057] <= 8'h86;
ROM_MEM[6058] <= 8'h07;
ROM_MEM[6059] <= 8'hA7;
ROM_MEM[6060] <= 8'h0C;
ROM_MEM[6061] <= 8'h86;
ROM_MEM[6062] <= 8'h18;
ROM_MEM[6063] <= 8'hA7;
ROM_MEM[6064] <= 8'h0D;
ROM_MEM[6065] <= 8'hEC;
ROM_MEM[6066] <= 8'h52;
ROM_MEM[6067] <= 8'hBD;
ROM_MEM[6068] <= 8'hCD;
ROM_MEM[6069] <= 8'h9C;
ROM_MEM[6070] <= 8'hED;
ROM_MEM[6071] <= 8'h06;
ROM_MEM[6072] <= 8'hE3;
ROM_MEM[6073] <= 8'h48;
ROM_MEM[6074] <= 8'hED;
ROM_MEM[6075] <= 8'h84;
ROM_MEM[6076] <= 8'hEC;
ROM_MEM[6077] <= 8'h5A;
ROM_MEM[6078] <= 8'hBD;
ROM_MEM[6079] <= 8'hCD;
ROM_MEM[6080] <= 8'h9C;
ROM_MEM[6081] <= 8'hED;
ROM_MEM[6082] <= 8'h08;
ROM_MEM[6083] <= 8'hE3;
ROM_MEM[6084] <= 8'h4A;
ROM_MEM[6085] <= 8'hED;
ROM_MEM[6086] <= 8'h02;
ROM_MEM[6087] <= 8'hEC;
ROM_MEM[6088] <= 8'h42;
ROM_MEM[6089] <= 8'hBD;
ROM_MEM[6090] <= 8'hCD;
ROM_MEM[6091] <= 8'h9C;
ROM_MEM[6092] <= 8'hED;
ROM_MEM[6093] <= 8'h0A;
ROM_MEM[6094] <= 8'hE3;
ROM_MEM[6095] <= 8'h4C;
ROM_MEM[6096] <= 8'hED;
ROM_MEM[6097] <= 8'h04;
ROM_MEM[6098] <= 8'hBD;
ROM_MEM[6099] <= 8'hB8;
ROM_MEM[6100] <= 8'h3F;
ROM_MEM[6101] <= 8'hBD;
ROM_MEM[6102] <= 8'hB9;
ROM_MEM[6103] <= 8'h48;
ROM_MEM[6104] <= 8'h86;
ROM_MEM[6105] <= 8'h08;
ROM_MEM[6106] <= 8'hA7;
ROM_MEM[6107] <= 8'h0C;
ROM_MEM[6108] <= 8'h86;
ROM_MEM[6109] <= 8'h10;
ROM_MEM[6110] <= 8'hA7;
ROM_MEM[6111] <= 8'h0D;
ROM_MEM[6112] <= 8'hEC;
ROM_MEM[6113] <= 8'h48;
ROM_MEM[6114] <= 8'hED;
ROM_MEM[6115] <= 8'h84;
ROM_MEM[6116] <= 8'hED;
ROM_MEM[6117] <= 8'h06;
ROM_MEM[6118] <= 8'hEC;
ROM_MEM[6119] <= 8'h4A;
ROM_MEM[6120] <= 8'hED;
ROM_MEM[6121] <= 8'h02;
ROM_MEM[6122] <= 8'hED;
ROM_MEM[6123] <= 8'h08;
ROM_MEM[6124] <= 8'hEC;
ROM_MEM[6125] <= 8'h4C;
ROM_MEM[6126] <= 8'hED;
ROM_MEM[6127] <= 8'h04;
ROM_MEM[6128] <= 8'hED;
ROM_MEM[6129] <= 8'h0A;
ROM_MEM[6130] <= 8'hA6;
ROM_MEM[6131] <= 8'h06;
ROM_MEM[6132] <= 8'hC6;
ROM_MEM[6133] <= 8'h80;
ROM_MEM[6134] <= 8'h58;
ROM_MEM[6135] <= 8'h49;
ROM_MEM[6136] <= 8'h28;
ROM_MEM[6137] <= 8'h04;
ROM_MEM[6138] <= 8'h46;
ROM_MEM[6139] <= 8'h56;
ROM_MEM[6140] <= 8'h20;
ROM_MEM[6141] <= 8'h1E;
ROM_MEM[6142] <= 8'h68;
ROM_MEM[6143] <= 8'h09;
ROM_MEM[6144] <= 8'h69;
ROM_MEM[6145] <= 8'h08;
ROM_MEM[6146] <= 8'h28;
ROM_MEM[6147] <= 8'h08;
ROM_MEM[6148] <= 8'h66;
ROM_MEM[6149] <= 8'h08;
ROM_MEM[6150] <= 8'h66;
ROM_MEM[6151] <= 8'h09;
ROM_MEM[6152] <= 8'h47;
ROM_MEM[6153] <= 8'h56;
ROM_MEM[6154] <= 8'h20;
ROM_MEM[6155] <= 8'h10;
ROM_MEM[6156] <= 8'h68;
ROM_MEM[6157] <= 8'h0B;
ROM_MEM[6158] <= 8'h69;
ROM_MEM[6159] <= 8'h0A;
ROM_MEM[6160] <= 8'h28;
ROM_MEM[6161] <= 8'hE4;
ROM_MEM[6162] <= 8'h66;
ROM_MEM[6163] <= 8'h0A;
ROM_MEM[6164] <= 8'h66;
ROM_MEM[6165] <= 8'h0B;
ROM_MEM[6166] <= 8'h67;
ROM_MEM[6167] <= 8'h08;
ROM_MEM[6168] <= 8'h67;
ROM_MEM[6169] <= 8'h09;
ROM_MEM[6170] <= 8'h47;
ROM_MEM[6171] <= 8'h56;
ROM_MEM[6172] <= 8'hA3;
ROM_MEM[6173] <= 8'h84;
ROM_MEM[6174] <= 8'hBD;
ROM_MEM[6175] <= 8'hCD;
ROM_MEM[6176] <= 8'hA0;
ROM_MEM[6177] <= 8'hF6;
ROM_MEM[6178] <= 8'h47;
ROM_MEM[6179] <= 8'h03;
ROM_MEM[6180] <= 8'hED;
ROM_MEM[6181] <= 8'h06;
ROM_MEM[6182] <= 8'hEC;
ROM_MEM[6183] <= 8'h08;
ROM_MEM[6184] <= 8'hA3;
ROM_MEM[6185] <= 8'h02;
ROM_MEM[6186] <= 8'hBD;
ROM_MEM[6187] <= 8'hCD;
ROM_MEM[6188] <= 8'hA0;
ROM_MEM[6189] <= 8'hF6;
ROM_MEM[6190] <= 8'h47;
ROM_MEM[6191] <= 8'h03;
ROM_MEM[6192] <= 8'hED;
ROM_MEM[6193] <= 8'h08;
ROM_MEM[6194] <= 8'hEC;
ROM_MEM[6195] <= 8'h0A;
ROM_MEM[6196] <= 8'hA3;
ROM_MEM[6197] <= 8'h04;
ROM_MEM[6198] <= 8'hBD;
ROM_MEM[6199] <= 8'hCD;
ROM_MEM[6200] <= 8'hA0;
ROM_MEM[6201] <= 8'hF6;
ROM_MEM[6202] <= 8'h47;
ROM_MEM[6203] <= 8'h03;
ROM_MEM[6204] <= 8'hED;
ROM_MEM[6205] <= 8'h0A;
ROM_MEM[6206] <= 8'h39;
ROM_MEM[6207] <= 8'hEC;
ROM_MEM[6208] <= 8'h56;
ROM_MEM[6209] <= 8'hE3;
ROM_MEM[6210] <= 8'h06;
ROM_MEM[6211] <= 8'hED;
ROM_MEM[6212] <= 8'h06;
ROM_MEM[6213] <= 8'hEC;
ROM_MEM[6214] <= 8'h5E;
ROM_MEM[6215] <= 8'hE3;
ROM_MEM[6216] <= 8'h08;
ROM_MEM[6217] <= 8'hED;
ROM_MEM[6218] <= 8'h08;
ROM_MEM[6219] <= 8'hEC;
ROM_MEM[6220] <= 8'h46;
ROM_MEM[6221] <= 8'hE3;
ROM_MEM[6222] <= 8'h0A;
ROM_MEM[6223] <= 8'hED;
ROM_MEM[6224] <= 8'h0A;
ROM_MEM[6225] <= 8'h39;
ROM_MEM[6226] <= 8'hCC;
ROM_MEM[6227] <= 8'h00;
ROM_MEM[6228] <= 8'h01;
ROM_MEM[6229] <= 8'hDD;
ROM_MEM[6230] <= 8'h01;
ROM_MEM[6231] <= 8'hCC;
ROM_MEM[6232] <= 8'h02;
ROM_MEM[6233] <= 8'h03;
ROM_MEM[6234] <= 8'hDD;
ROM_MEM[6235] <= 8'h03;
ROM_MEM[6236] <= 8'h20;
ROM_MEM[6237] <= 8'h0A;
ROM_MEM[6238] <= 8'hCC;
ROM_MEM[6239] <= 8'h03;
ROM_MEM[6240] <= 8'h04;
ROM_MEM[6241] <= 8'hDD;
ROM_MEM[6242] <= 8'h01;
ROM_MEM[6243] <= 8'hCC;
ROM_MEM[6244] <= 8'h05;
ROM_MEM[6245] <= 8'h02;
ROM_MEM[6246] <= 8'hDD;
ROM_MEM[6247] <= 8'h03;
ROM_MEM[6248] <= 8'hBD;
ROM_MEM[6249] <= 8'hB9;
ROM_MEM[6250] <= 8'h48;
ROM_MEM[6251] <= 8'h96;
ROM_MEM[6252] <= 8'h01;
ROM_MEM[6253] <= 8'hA7;
ROM_MEM[6254] <= 8'h0C;
ROM_MEM[6255] <= 8'h86;
ROM_MEM[6256] <= 8'h20;
ROM_MEM[6257] <= 8'hA7;
ROM_MEM[6258] <= 8'h0D;
ROM_MEM[6259] <= 8'hFC;
ROM_MEM[6260] <= 8'h50;
ROM_MEM[6261] <= 8'h18;
ROM_MEM[6262] <= 8'hED;
ROM_MEM[6263] <= 8'h84;
ROM_MEM[6264] <= 8'hFC;
ROM_MEM[6265] <= 8'h50;
ROM_MEM[6266] <= 8'h1A;
ROM_MEM[6267] <= 8'h8B;
ROM_MEM[6268] <= 8'hFE;
ROM_MEM[6269] <= 8'hED;
ROM_MEM[6270] <= 8'h02;
ROM_MEM[6271] <= 8'hFC;
ROM_MEM[6272] <= 8'h50;
ROM_MEM[6273] <= 8'h1C;
ROM_MEM[6274] <= 8'hED;
ROM_MEM[6275] <= 8'h04;
ROM_MEM[6276] <= 8'hFC;
ROM_MEM[6277] <= 8'h50;
ROM_MEM[6278] <= 8'h98;
ROM_MEM[6279] <= 8'h8B;
ROM_MEM[6280] <= 8'h7F;
ROM_MEM[6281] <= 8'hB3;
ROM_MEM[6282] <= 8'h50;
ROM_MEM[6283] <= 8'h18;
ROM_MEM[6284] <= 8'hBD;
ROM_MEM[6285] <= 8'hCD;
ROM_MEM[6286] <= 8'h9E;
ROM_MEM[6287] <= 8'hF6;
ROM_MEM[6288] <= 8'h47;
ROM_MEM[6289] <= 8'h03;
ROM_MEM[6290] <= 8'hED;
ROM_MEM[6291] <= 8'h06;
ROM_MEM[6292] <= 8'hFC;
ROM_MEM[6293] <= 8'h50;
ROM_MEM[6294] <= 8'h9A;
ROM_MEM[6295] <= 8'h8B;
ROM_MEM[6296] <= 8'hC1;
ROM_MEM[6297] <= 8'hB3;
ROM_MEM[6298] <= 8'h50;
ROM_MEM[6299] <= 8'h1A;
ROM_MEM[6300] <= 8'hBD;
ROM_MEM[6301] <= 8'hCD;
ROM_MEM[6302] <= 8'h9E;
ROM_MEM[6303] <= 8'hF6;
ROM_MEM[6304] <= 8'h47;
ROM_MEM[6305] <= 8'h03;
ROM_MEM[6306] <= 8'hED;
ROM_MEM[6307] <= 8'h08;
ROM_MEM[6308] <= 8'h96;
ROM_MEM[6309] <= 8'h04;
ROM_MEM[6310] <= 8'hF6;
ROM_MEM[6311] <= 8'h47;
ROM_MEM[6312] <= 8'h03;
ROM_MEM[6313] <= 8'hBD;
ROM_MEM[6314] <= 8'hCD;
ROM_MEM[6315] <= 8'hB5;
ROM_MEM[6316] <= 8'hED;
ROM_MEM[6317] <= 8'h0A;
ROM_MEM[6318] <= 8'hBD;
ROM_MEM[6319] <= 8'hB9;
ROM_MEM[6320] <= 8'h48;
ROM_MEM[6321] <= 8'h96;
ROM_MEM[6322] <= 8'h02;
ROM_MEM[6323] <= 8'hA7;
ROM_MEM[6324] <= 8'h0C;
ROM_MEM[6325] <= 8'h86;
ROM_MEM[6326] <= 8'h20;
ROM_MEM[6327] <= 8'hA7;
ROM_MEM[6328] <= 8'h0D;
ROM_MEM[6329] <= 8'hFC;
ROM_MEM[6330] <= 8'h50;
ROM_MEM[6331] <= 8'h18;
ROM_MEM[6332] <= 8'h8B;
ROM_MEM[6333] <= 8'h02;
ROM_MEM[6334] <= 8'hED;
ROM_MEM[6335] <= 8'h84;
ROM_MEM[6336] <= 8'hFC;
ROM_MEM[6337] <= 8'h50;
ROM_MEM[6338] <= 8'h1A;
ROM_MEM[6339] <= 8'hED;
ROM_MEM[6340] <= 8'h02;
ROM_MEM[6341] <= 8'hFC;
ROM_MEM[6342] <= 8'h50;
ROM_MEM[6343] <= 8'h1C;
ROM_MEM[6344] <= 8'hED;
ROM_MEM[6345] <= 8'h04;
ROM_MEM[6346] <= 8'hFC;
ROM_MEM[6347] <= 8'h50;
ROM_MEM[6348] <= 8'h98;
ROM_MEM[6349] <= 8'h8B;
ROM_MEM[6350] <= 8'h7F;
ROM_MEM[6351] <= 8'hB3;
ROM_MEM[6352] <= 8'h50;
ROM_MEM[6353] <= 8'h18;
ROM_MEM[6354] <= 8'hBD;
ROM_MEM[6355] <= 8'hCD;
ROM_MEM[6356] <= 8'h9E;
ROM_MEM[6357] <= 8'hF6;
ROM_MEM[6358] <= 8'h47;
ROM_MEM[6359] <= 8'h03;
ROM_MEM[6360] <= 8'hED;
ROM_MEM[6361] <= 8'h06;
ROM_MEM[6362] <= 8'hFC;
ROM_MEM[6363] <= 8'h50;
ROM_MEM[6364] <= 8'h9A;
ROM_MEM[6365] <= 8'hB3;
ROM_MEM[6366] <= 8'h50;
ROM_MEM[6367] <= 8'h1A;
ROM_MEM[6368] <= 8'hBD;
ROM_MEM[6369] <= 8'hCD;
ROM_MEM[6370] <= 8'h9E;
ROM_MEM[6371] <= 8'hF6;
ROM_MEM[6372] <= 8'h47;
ROM_MEM[6373] <= 8'h03;
ROM_MEM[6374] <= 8'hED;
ROM_MEM[6375] <= 8'h08;
ROM_MEM[6376] <= 8'h96;
ROM_MEM[6377] <= 8'h04;
ROM_MEM[6378] <= 8'hF6;
ROM_MEM[6379] <= 8'h47;
ROM_MEM[6380] <= 8'h03;
ROM_MEM[6381] <= 8'hBD;
ROM_MEM[6382] <= 8'hCD;
ROM_MEM[6383] <= 8'hB5;
ROM_MEM[6384] <= 8'hED;
ROM_MEM[6385] <= 8'h0A;
ROM_MEM[6386] <= 8'hBD;
ROM_MEM[6387] <= 8'hB9;
ROM_MEM[6388] <= 8'h48;
ROM_MEM[6389] <= 8'h96;
ROM_MEM[6390] <= 8'h03;
ROM_MEM[6391] <= 8'hA7;
ROM_MEM[6392] <= 8'h0C;
ROM_MEM[6393] <= 8'h86;
ROM_MEM[6394] <= 8'h20;
ROM_MEM[6395] <= 8'hA7;
ROM_MEM[6396] <= 8'h0D;
ROM_MEM[6397] <= 8'hFC;
ROM_MEM[6398] <= 8'h50;
ROM_MEM[6399] <= 8'h18;
ROM_MEM[6400] <= 8'hED;
ROM_MEM[6401] <= 8'h84;
ROM_MEM[6402] <= 8'hFC;
ROM_MEM[6403] <= 8'h50;
ROM_MEM[6404] <= 8'h1A;
ROM_MEM[6405] <= 8'h8B;
ROM_MEM[6406] <= 8'h02;
ROM_MEM[6407] <= 8'hED;
ROM_MEM[6408] <= 8'h02;
ROM_MEM[6409] <= 8'hFC;
ROM_MEM[6410] <= 8'h50;
ROM_MEM[6411] <= 8'h1C;
ROM_MEM[6412] <= 8'hED;
ROM_MEM[6413] <= 8'h04;
ROM_MEM[6414] <= 8'hFC;
ROM_MEM[6415] <= 8'h50;
ROM_MEM[6416] <= 8'h98;
ROM_MEM[6417] <= 8'h8B;
ROM_MEM[6418] <= 8'h7F;
ROM_MEM[6419] <= 8'hB3;
ROM_MEM[6420] <= 8'h50;
ROM_MEM[6421] <= 8'h18;
ROM_MEM[6422] <= 8'hBD;
ROM_MEM[6423] <= 8'hCD;
ROM_MEM[6424] <= 8'h9E;
ROM_MEM[6425] <= 8'hF6;
ROM_MEM[6426] <= 8'h47;
ROM_MEM[6427] <= 8'h03;
ROM_MEM[6428] <= 8'hED;
ROM_MEM[6429] <= 8'h06;
ROM_MEM[6430] <= 8'hFC;
ROM_MEM[6431] <= 8'h50;
ROM_MEM[6432] <= 8'h9A;
ROM_MEM[6433] <= 8'h8B;
ROM_MEM[6434] <= 8'h3F;
ROM_MEM[6435] <= 8'hB3;
ROM_MEM[6436] <= 8'h50;
ROM_MEM[6437] <= 8'h1A;
ROM_MEM[6438] <= 8'hBD;
ROM_MEM[6439] <= 8'hCD;
ROM_MEM[6440] <= 8'h9E;
ROM_MEM[6441] <= 8'hF6;
ROM_MEM[6442] <= 8'h47;
ROM_MEM[6443] <= 8'h03;
ROM_MEM[6444] <= 8'hED;
ROM_MEM[6445] <= 8'h08;
ROM_MEM[6446] <= 8'h96;
ROM_MEM[6447] <= 8'h04;
ROM_MEM[6448] <= 8'hF6;
ROM_MEM[6449] <= 8'h47;
ROM_MEM[6450] <= 8'h03;
ROM_MEM[6451] <= 8'hBD;
ROM_MEM[6452] <= 8'hCD;
ROM_MEM[6453] <= 8'hB5;
ROM_MEM[6454] <= 8'hED;
ROM_MEM[6455] <= 8'h0A;
ROM_MEM[6456] <= 8'h39;
ROM_MEM[6457] <= 8'h8E;
ROM_MEM[6458] <= 8'h49;
ROM_MEM[6459] <= 8'hE2;
ROM_MEM[6460] <= 8'h86;
ROM_MEM[6461] <= 8'h00;
ROM_MEM[6462] <= 8'hA7;
ROM_MEM[6463] <= 8'h0D;
ROM_MEM[6464] <= 8'h30;
ROM_MEM[6465] <= 8'h0E;
ROM_MEM[6466] <= 8'h8C;
ROM_MEM[6467] <= 8'h4A;
ROM_MEM[6468] <= 8'h52;
ROM_MEM[6469] <= 8'h25;
ROM_MEM[6470] <= 8'hF5;
ROM_MEM[6471] <= 8'h39;
ROM_MEM[6472] <= 8'hD6;
ROM_MEM[6473] <= 8'hA2;
ROM_MEM[6474] <= 8'h5C;
ROM_MEM[6475] <= 8'hC1;
ROM_MEM[6476] <= 8'h08;
ROM_MEM[6477] <= 8'h25;
ROM_MEM[6478] <= 8'h02;
ROM_MEM[6479] <= 8'hC6;
ROM_MEM[6480] <= 8'h00;
ROM_MEM[6481] <= 8'hD7;
ROM_MEM[6482] <= 8'hA2;
ROM_MEM[6483] <= 8'h86;
ROM_MEM[6484] <= 8'h0E;
ROM_MEM[6485] <= 8'h3D;
ROM_MEM[6486] <= 8'h8E;
ROM_MEM[6487] <= 8'h49;
ROM_MEM[6488] <= 8'hE2;
ROM_MEM[6489] <= 8'h30;
ROM_MEM[6490] <= 8'h8B;
ROM_MEM[6491] <= 8'h39;
ROM_MEM[6492] <= 8'hCC;
ROM_MEM[6493] <= 8'h14;
ROM_MEM[6494] <= 8'hBD;
ROM_MEM[6495] <= 8'hFD;
ROM_MEM[6496] <= 8'h50;
ROM_MEM[6497] <= 8'h22;
ROM_MEM[6498] <= 8'hCC;
ROM_MEM[6499] <= 8'h3C;
ROM_MEM[6500] <= 8'h8C;
ROM_MEM[6501] <= 8'hFD;
ROM_MEM[6502] <= 8'h50;
ROM_MEM[6503] <= 8'h24;
ROM_MEM[6504] <= 8'hCC;
ROM_MEM[6505] <= 8'h00;
ROM_MEM[6506] <= 8'h18;
ROM_MEM[6507] <= 8'hFD;
ROM_MEM[6508] <= 8'h47;
ROM_MEM[6509] <= 8'h01;
ROM_MEM[6510] <= 8'h86;
ROM_MEM[6511] <= 8'h00;
ROM_MEM[6512] <= 8'hBD;
ROM_MEM[6513] <= 8'hCD;
ROM_MEM[6514] <= 8'hBA;
ROM_MEM[6515] <= 8'hCC;
ROM_MEM[6516] <= 8'h05;
ROM_MEM[6517] <= 8'h90;
ROM_MEM[6518] <= 8'hFD;
ROM_MEM[6519] <= 8'h50;
ROM_MEM[6520] <= 8'h22;
ROM_MEM[6521] <= 8'hCC;
ROM_MEM[6522] <= 8'h3F;
ROM_MEM[6523] <= 8'hC2;
ROM_MEM[6524] <= 8'hFD;
ROM_MEM[6525] <= 8'h50;
ROM_MEM[6526] <= 8'h24;
ROM_MEM[6527] <= 8'hCC;
ROM_MEM[6528] <= 8'h00;
ROM_MEM[6529] <= 8'h18;
ROM_MEM[6530] <= 8'hFD;
ROM_MEM[6531] <= 8'h47;
ROM_MEM[6532] <= 8'h01;
ROM_MEM[6533] <= 8'h86;
ROM_MEM[6534] <= 8'h0E;
ROM_MEM[6535] <= 8'hBD;
ROM_MEM[6536] <= 8'hCD;
ROM_MEM[6537] <= 8'hBA;
ROM_MEM[6538] <= 8'h39;
ROM_MEM[6539] <= 8'h8E;
ROM_MEM[6540] <= 8'h49;
ROM_MEM[6541] <= 8'hE2;
ROM_MEM[6542] <= 8'hA6;
ROM_MEM[6543] <= 8'h0D;
ROM_MEM[6544] <= 8'h27;
ROM_MEM[6545] <= 8'h0F;
ROM_MEM[6546] <= 8'h6A;
ROM_MEM[6547] <= 8'h0D;
ROM_MEM[6548] <= 8'hE6;
ROM_MEM[6549] <= 8'h0C;
ROM_MEM[6550] <= 8'hC1;
ROM_MEM[6551] <= 8'h09;
ROM_MEM[6552] <= 8'h25;
ROM_MEM[6553] <= 8'h01;
ROM_MEM[6554] <= 8'h3F;
ROM_MEM[6555] <= 8'hCE;
ROM_MEM[6556] <= 8'hB7;
ROM_MEM[6557] <= 8'h48;
ROM_MEM[6558] <= 8'h58;
ROM_MEM[6559] <= 8'hAD;
ROM_MEM[6560] <= 8'hD5;
ROM_MEM[6561] <= 8'h30;
ROM_MEM[6562] <= 8'h0E;
ROM_MEM[6563] <= 8'h8C;
ROM_MEM[6564] <= 8'h4A;
ROM_MEM[6565] <= 8'h52;
ROM_MEM[6566] <= 8'h25;
ROM_MEM[6567] <= 8'hE6;
ROM_MEM[6568] <= 8'h8E;
ROM_MEM[6569] <= 8'h49;
ROM_MEM[6570] <= 8'hE2;
ROM_MEM[6571] <= 8'hA6;
ROM_MEM[6572] <= 8'h0D;
ROM_MEM[6573] <= 8'h27;
ROM_MEM[6574] <= 8'h03;
ROM_MEM[6575] <= 8'h7E;
ROM_MEM[6576] <= 8'hB9;
ROM_MEM[6577] <= 8'h5C;
ROM_MEM[6578] <= 8'h30;
ROM_MEM[6579] <= 8'h0E;
ROM_MEM[6580] <= 8'h8C;
ROM_MEM[6581] <= 8'h4A;
ROM_MEM[6582] <= 8'h52;
ROM_MEM[6583] <= 8'h25;
ROM_MEM[6584] <= 8'hF2;
ROM_MEM[6585] <= 8'hCE;
ROM_MEM[6586] <= 8'h50;
ROM_MEM[6587] <= 8'hD0;
ROM_MEM[6588] <= 8'hBD;
ROM_MEM[6589] <= 8'hCD;
ROM_MEM[6590] <= 8'hC3;
ROM_MEM[6591] <= 8'h39;
ROM_MEM[6592] <= 8'hEC;
ROM_MEM[6593] <= 8'h06;
ROM_MEM[6594] <= 8'hE3;
ROM_MEM[6595] <= 8'h84;
ROM_MEM[6596] <= 8'hED;
ROM_MEM[6597] <= 8'h84;
ROM_MEM[6598] <= 8'hCC;
ROM_MEM[6599] <= 8'h00;
ROM_MEM[6600] <= 8'h00;
ROM_MEM[6601] <= 8'hA3;
ROM_MEM[6602] <= 8'h06;
ROM_MEM[6603] <= 8'hBD;
ROM_MEM[6604] <= 8'hCD;
ROM_MEM[6605] <= 8'h9E;
ROM_MEM[6606] <= 8'hE3;
ROM_MEM[6607] <= 8'h06;
ROM_MEM[6608] <= 8'hED;
ROM_MEM[6609] <= 8'h06;
ROM_MEM[6610] <= 8'hEC;
ROM_MEM[6611] <= 8'h08;
ROM_MEM[6612] <= 8'hE3;
ROM_MEM[6613] <= 8'h02;
ROM_MEM[6614] <= 8'hED;
ROM_MEM[6615] <= 8'h02;
ROM_MEM[6616] <= 8'hCC;
ROM_MEM[6617] <= 8'h00;
ROM_MEM[6618] <= 8'h00;
ROM_MEM[6619] <= 8'hA3;
ROM_MEM[6620] <= 8'h08;
ROM_MEM[6621] <= 8'hBD;
ROM_MEM[6622] <= 8'hCD;
ROM_MEM[6623] <= 8'h9E;
ROM_MEM[6624] <= 8'hE3;
ROM_MEM[6625] <= 8'h08;
ROM_MEM[6626] <= 8'hED;
ROM_MEM[6627] <= 8'h08;
ROM_MEM[6628] <= 8'hEC;
ROM_MEM[6629] <= 8'h04;
ROM_MEM[6630] <= 8'hE3;
ROM_MEM[6631] <= 8'h0A;
ROM_MEM[6632] <= 8'h29;
ROM_MEM[6633] <= 8'h07;
ROM_MEM[6634] <= 8'h2C;
ROM_MEM[6635] <= 8'h03;
ROM_MEM[6636] <= 8'hCC;
ROM_MEM[6637] <= 8'h00;
ROM_MEM[6638] <= 8'h00;
ROM_MEM[6639] <= 8'hED;
ROM_MEM[6640] <= 8'h04;
ROM_MEM[6641] <= 8'hEC;
ROM_MEM[6642] <= 8'h0A;
ROM_MEM[6643] <= 8'h83;
ROM_MEM[6644] <= 8'h00;
ROM_MEM[6645] <= 8'hC8;
ROM_MEM[6646] <= 8'hED;
ROM_MEM[6647] <= 8'h0A;
ROM_MEM[6648] <= 8'h39;
ROM_MEM[6649] <= 8'hEC;
ROM_MEM[6650] <= 8'h06;
ROM_MEM[6651] <= 8'hE3;
ROM_MEM[6652] <= 8'h84;
ROM_MEM[6653] <= 8'h29;
ROM_MEM[6654] <= 8'h02;
ROM_MEM[6655] <= 8'hED;
ROM_MEM[6656] <= 8'h84;
ROM_MEM[6657] <= 8'hEC;
ROM_MEM[6658] <= 8'h08;
ROM_MEM[6659] <= 8'hE3;
ROM_MEM[6660] <= 8'h02;
ROM_MEM[6661] <= 8'h29;
ROM_MEM[6662] <= 8'h02;
ROM_MEM[6663] <= 8'hED;
ROM_MEM[6664] <= 8'h02;
ROM_MEM[6665] <= 8'hEC;
ROM_MEM[6666] <= 8'h0A;
ROM_MEM[6667] <= 8'hE3;
ROM_MEM[6668] <= 8'h04;
ROM_MEM[6669] <= 8'h29;
ROM_MEM[6670] <= 8'h02;
ROM_MEM[6671] <= 8'hED;
ROM_MEM[6672] <= 8'h04;
ROM_MEM[6673] <= 8'h39;
ROM_MEM[6674] <= 8'h86;
ROM_MEM[6675] <= 8'h18;
ROM_MEM[6676] <= 8'hBD;
ROM_MEM[6677] <= 8'hCE;
ROM_MEM[6678] <= 8'h18;
ROM_MEM[6679] <= 8'h86;
ROM_MEM[6680] <= 8'h40;
ROM_MEM[6681] <= 8'hBD;
ROM_MEM[6682] <= 8'hCD;
ROM_MEM[6683] <= 8'hBA;
ROM_MEM[6684] <= 8'h8E;
ROM_MEM[6685] <= 8'h49;
ROM_MEM[6686] <= 8'hE2;
ROM_MEM[6687] <= 8'h9F;
ROM_MEM[6688] <= 8'h64;
ROM_MEM[6689] <= 8'hA6;
ROM_MEM[6690] <= 8'h0D;
ROM_MEM[6691] <= 8'h27;
ROM_MEM[6692] <= 8'h03;
ROM_MEM[6693] <= 8'hBD;
ROM_MEM[6694] <= 8'hBA;
ROM_MEM[6695] <= 8'h32;
ROM_MEM[6696] <= 8'h9E;
ROM_MEM[6697] <= 8'h64;
ROM_MEM[6698] <= 8'h30;
ROM_MEM[6699] <= 8'h0E;
ROM_MEM[6700] <= 8'h8C;
ROM_MEM[6701] <= 8'h4A;
ROM_MEM[6702] <= 8'h52;
ROM_MEM[6703] <= 8'h25;
ROM_MEM[6704] <= 8'hEE;
ROM_MEM[6705] <= 8'h39;
ROM_MEM[6706] <= 8'hEC;
ROM_MEM[6707] <= 8'h84;
ROM_MEM[6708] <= 8'hFD;
ROM_MEM[6709] <= 8'h50;
ROM_MEM[6710] <= 8'h78;
ROM_MEM[6711] <= 8'hEC;
ROM_MEM[6712] <= 8'h02;
ROM_MEM[6713] <= 8'hFD;
ROM_MEM[6714] <= 8'h50;
ROM_MEM[6715] <= 8'h7A;
ROM_MEM[6716] <= 8'hEC;
ROM_MEM[6717] <= 8'h04;
ROM_MEM[6718] <= 8'hFD;
ROM_MEM[6719] <= 8'h50;
ROM_MEM[6720] <= 8'h7C;
ROM_MEM[6721] <= 8'hCC;
ROM_MEM[6722] <= 8'h00;
ROM_MEM[6723] <= 8'h0F;
ROM_MEM[6724] <= 8'hFD;
ROM_MEM[6725] <= 8'h47;
ROM_MEM[6726] <= 8'h01;
ROM_MEM[6727] <= 8'h86;
ROM_MEM[6728] <= 8'h67;
ROM_MEM[6729] <= 8'hBD;
ROM_MEM[6730] <= 8'hCD;
ROM_MEM[6731] <= 8'hBA;
ROM_MEM[6732] <= 8'hFC;
ROM_MEM[6733] <= 8'h50;
ROM_MEM[6734] <= 8'h00;
ROM_MEM[6735] <= 8'h2B;
ROM_MEM[6736] <= 8'h4C;
ROM_MEM[6737] <= 8'hFD;
ROM_MEM[6738] <= 8'h50;
ROM_MEM[6739] <= 8'h18;
ROM_MEM[6740] <= 8'hFD;
ROM_MEM[6741] <= 8'h47;
ROM_MEM[6742] <= 8'h04;
ROM_MEM[6743] <= 8'hFC;
ROM_MEM[6744] <= 8'h50;
ROM_MEM[6745] <= 8'h02;
ROM_MEM[6746] <= 8'hFD;
ROM_MEM[6747] <= 8'h50;
ROM_MEM[6748] <= 8'h1A;
ROM_MEM[6749] <= 8'h2A;
ROM_MEM[6750] <= 8'h04;
ROM_MEM[6751] <= 8'h43;
ROM_MEM[6752] <= 8'h50;
ROM_MEM[6753] <= 8'h82;
ROM_MEM[6754] <= 8'hFF;
ROM_MEM[6755] <= 8'hB3;
ROM_MEM[6756] <= 8'h50;
ROM_MEM[6757] <= 8'h18;
ROM_MEM[6758] <= 8'h2C;
ROM_MEM[6759] <= 8'h35;
ROM_MEM[6760] <= 8'hFC;
ROM_MEM[6761] <= 8'h50;
ROM_MEM[6762] <= 8'h04;
ROM_MEM[6763] <= 8'hFD;
ROM_MEM[6764] <= 8'h50;
ROM_MEM[6765] <= 8'h1C;
ROM_MEM[6766] <= 8'h2A;
ROM_MEM[6767] <= 8'h04;
ROM_MEM[6768] <= 8'h43;
ROM_MEM[6769] <= 8'h50;
ROM_MEM[6770] <= 8'h82;
ROM_MEM[6771] <= 8'hFF;
ROM_MEM[6772] <= 8'h44;
ROM_MEM[6773] <= 8'h56;
ROM_MEM[6774] <= 8'hB3;
ROM_MEM[6775] <= 8'h50;
ROM_MEM[6776] <= 8'h18;
ROM_MEM[6777] <= 8'h2C;
ROM_MEM[6778] <= 8'h22;
ROM_MEM[6779] <= 8'hE6;
ROM_MEM[6780] <= 8'h0C;
ROM_MEM[6781] <= 8'hC1;
ROM_MEM[6782] <= 8'h09;
ROM_MEM[6783] <= 8'h25;
ROM_MEM[6784] <= 8'h01;
ROM_MEM[6785] <= 8'h3F;
ROM_MEM[6786] <= 8'hCE;
ROM_MEM[6787] <= 8'hB7;
ROM_MEM[6788] <= 8'h5A;
ROM_MEM[6789] <= 8'h58;
ROM_MEM[6790] <= 8'hAD;
ROM_MEM[6791] <= 8'hD5;
ROM_MEM[6792] <= 8'hBD;
ROM_MEM[6793] <= 8'hCC;
ROM_MEM[6794] <= 8'hD8;
ROM_MEM[6795] <= 8'hBD;
ROM_MEM[6796] <= 8'hCD;
ROM_MEM[6797] <= 8'h20;
ROM_MEM[6798] <= 8'hBD;
ROM_MEM[6799] <= 8'hCD;
ROM_MEM[6800] <= 8'h2C;
ROM_MEM[6801] <= 8'hCC;
ROM_MEM[6802] <= 8'h72;
ROM_MEM[6803] <= 8'h00;
ROM_MEM[6804] <= 8'hED;
ROM_MEM[6805] <= 8'hA1;
ROM_MEM[6806] <= 8'hCC;
ROM_MEM[6807] <= 8'h80;
ROM_MEM[6808] <= 8'h40;
ROM_MEM[6809] <= 8'hED;
ROM_MEM[6810] <= 8'hA1;
ROM_MEM[6811] <= 8'h20;
ROM_MEM[6812] <= 8'h02;
ROM_MEM[6813] <= 8'h6F;
ROM_MEM[6814] <= 8'h0D;
ROM_MEM[6815] <= 8'h39;
ROM_MEM[6816] <= 8'h86;
ROM_MEM[6817] <= 8'h14;
ROM_MEM[6818] <= 8'h20;
ROM_MEM[6819] <= 8'h1A;
ROM_MEM[6820] <= 8'h86;
ROM_MEM[6821] <= 8'h15;
ROM_MEM[6822] <= 8'h20;
ROM_MEM[6823] <= 8'h16;
ROM_MEM[6824] <= 8'h86;
ROM_MEM[6825] <= 8'h16;
ROM_MEM[6826] <= 8'h20;
ROM_MEM[6827] <= 8'h12;
ROM_MEM[6828] <= 8'h86;
ROM_MEM[6829] <= 8'h11;
ROM_MEM[6830] <= 8'h20;
ROM_MEM[6831] <= 8'h08;
ROM_MEM[6832] <= 8'h86;
ROM_MEM[6833] <= 8'h12;
ROM_MEM[6834] <= 8'h20;
ROM_MEM[6835] <= 8'h04;
ROM_MEM[6836] <= 8'h86;
ROM_MEM[6837] <= 8'h13;
ROM_MEM[6838] <= 8'h20;
ROM_MEM[6839] <= 8'h00;
ROM_MEM[6840] <= 8'h97;
ROM_MEM[6841] <= 8'hDC;
ROM_MEM[6842] <= 8'h86;
ROM_MEM[6843] <= 8'h67;
ROM_MEM[6844] <= 8'h20;
ROM_MEM[6845] <= 8'h04;
ROM_MEM[6846] <= 8'h97;
ROM_MEM[6847] <= 8'hDC;
ROM_MEM[6848] <= 8'h86;
ROM_MEM[6849] <= 8'h64;
ROM_MEM[6850] <= 8'hE6;
ROM_MEM[6851] <= 8'h0D;
ROM_MEM[6852] <= 8'hC1;
ROM_MEM[6853] <= 8'h07;
ROM_MEM[6854] <= 8'h22;
ROM_MEM[6855] <= 8'h06;
ROM_MEM[6856] <= 8'h58;
ROM_MEM[6857] <= 8'h58;
ROM_MEM[6858] <= 8'h58;
ROM_MEM[6859] <= 8'h58;
ROM_MEM[6860] <= 8'h20;
ROM_MEM[6861] <= 8'h02;
ROM_MEM[6862] <= 8'hC6;
ROM_MEM[6863] <= 8'h80;
ROM_MEM[6864] <= 8'hED;
ROM_MEM[6865] <= 8'hA1;
ROM_MEM[6866] <= 8'hEC;
ROM_MEM[6867] <= 8'h84;
ROM_MEM[6868] <= 8'hFD;
ROM_MEM[6869] <= 8'h50;
ROM_MEM[6870] <= 8'h78;
ROM_MEM[6871] <= 8'hEC;
ROM_MEM[6872] <= 8'h02;
ROM_MEM[6873] <= 8'hFD;
ROM_MEM[6874] <= 8'h50;
ROM_MEM[6875] <= 8'h7A;
ROM_MEM[6876] <= 8'hCC;
ROM_MEM[6877] <= 8'h00;
ROM_MEM[6878] <= 8'h00;
ROM_MEM[6879] <= 8'hFD;
ROM_MEM[6880] <= 8'h50;
ROM_MEM[6881] <= 8'h7C;
ROM_MEM[6882] <= 8'hCC;
ROM_MEM[6883] <= 8'h00;
ROM_MEM[6884] <= 8'h0F;
ROM_MEM[6885] <= 8'hFD;
ROM_MEM[6886] <= 8'h47;
ROM_MEM[6887] <= 8'h01;
ROM_MEM[6888] <= 8'hFC;
ROM_MEM[6889] <= 8'h50;
ROM_MEM[6890] <= 8'h1C;
ROM_MEM[6891] <= 8'h34;
ROM_MEM[6892] <= 8'h56;
ROM_MEM[6893] <= 8'hFE;
ROM_MEM[6894] <= 8'h50;
ROM_MEM[6895] <= 8'h1A;
ROM_MEM[6896] <= 8'hBE;
ROM_MEM[6897] <= 8'h50;
ROM_MEM[6898] <= 8'h18;
ROM_MEM[6899] <= 8'h86;
ROM_MEM[6900] <= 8'h67;
ROM_MEM[6901] <= 8'hBD;
ROM_MEM[6902] <= 8'hCD;
ROM_MEM[6903] <= 8'hBA;
ROM_MEM[6904] <= 8'hBF;
ROM_MEM[6905] <= 8'h50;
ROM_MEM[6906] <= 8'h18;
ROM_MEM[6907] <= 8'hFF;
ROM_MEM[6908] <= 8'h50;
ROM_MEM[6909] <= 8'h1A;
ROM_MEM[6910] <= 8'h35;
ROM_MEM[6911] <= 8'h56;
ROM_MEM[6912] <= 8'hFD;
ROM_MEM[6913] <= 8'h50;
ROM_MEM[6914] <= 8'h1C;
ROM_MEM[6915] <= 8'hFC;
ROM_MEM[6916] <= 8'h50;
ROM_MEM[6917] <= 8'h00;
ROM_MEM[6918] <= 8'hFD;
ROM_MEM[6919] <= 8'h47;
ROM_MEM[6920] <= 8'h04;
ROM_MEM[6921] <= 8'hBD;
ROM_MEM[6922] <= 8'hCC;
ROM_MEM[6923] <= 8'hF0;
ROM_MEM[6924] <= 8'h86;
ROM_MEM[6925] <= 8'h72;
ROM_MEM[6926] <= 8'hF6;
ROM_MEM[6927] <= 8'h50;
ROM_MEM[6928] <= 8'h18;
ROM_MEM[6929] <= 8'h58;
ROM_MEM[6930] <= 8'h58;
ROM_MEM[6931] <= 8'hED;
ROM_MEM[6932] <= 8'hA1;
ROM_MEM[6933] <= 8'h39;
ROM_MEM[6934] <= 8'hC6;
ROM_MEM[6935] <= 8'h03;
ROM_MEM[6936] <= 8'h20;
ROM_MEM[6937] <= 8'h08;
ROM_MEM[6938] <= 8'hC6;
ROM_MEM[6939] <= 8'h01;
ROM_MEM[6940] <= 8'h20;
ROM_MEM[6941] <= 8'h04;
ROM_MEM[6942] <= 8'hC6;
ROM_MEM[6943] <= 8'h02;
ROM_MEM[6944] <= 8'h20;
ROM_MEM[6945] <= 8'h00;
ROM_MEM[6946] <= 8'hD7;
ROM_MEM[6947] <= 8'hDC;
ROM_MEM[6948] <= 8'hE6;
ROM_MEM[6949] <= 8'h0D;
ROM_MEM[6950] <= 8'hC1;
ROM_MEM[6951] <= 8'h1F;
ROM_MEM[6952] <= 8'h23;
ROM_MEM[6953] <= 8'h05;
ROM_MEM[6954] <= 8'hCC;
ROM_MEM[6955] <= 8'hA0;
ROM_MEM[6956] <= 8'h18;
ROM_MEM[6957] <= 8'h20;
ROM_MEM[6958] <= 8'h06;
ROM_MEM[6959] <= 8'hCE;
ROM_MEM[6960] <= 8'hBB;
ROM_MEM[6961] <= 8'h3B;
ROM_MEM[6962] <= 8'h58;
ROM_MEM[6963] <= 8'hEC;
ROM_MEM[6964] <= 8'hC5;
ROM_MEM[6965] <= 8'hED;
ROM_MEM[6966] <= 8'hA1;
ROM_MEM[6967] <= 8'hBD;
ROM_MEM[6968] <= 8'hCC;
ROM_MEM[6969] <= 8'hF0;
ROM_MEM[6970] <= 8'h39;
ROM_MEM[6971] <= 8'h62;
ROM_MEM[6972] <= 8'h30;
ROM_MEM[6973] <= 8'h62;
ROM_MEM[6974] <= 8'h30;
ROM_MEM[6975] <= 8'h62;
ROM_MEM[6976] <= 8'h40;
ROM_MEM[6977] <= 8'h62;
ROM_MEM[6978] <= 8'h40;
ROM_MEM[6979] <= 8'h62;
ROM_MEM[6980] <= 8'h50;
ROM_MEM[6981] <= 8'h62;
ROM_MEM[6982] <= 8'h50;
ROM_MEM[6983] <= 8'h62;
ROM_MEM[6984] <= 8'h60;
ROM_MEM[6985] <= 8'h62;
ROM_MEM[6986] <= 8'h60;
ROM_MEM[6987] <= 8'h62;
ROM_MEM[6988] <= 8'h70;
ROM_MEM[6989] <= 8'h62;
ROM_MEM[6990] <= 8'h70;
ROM_MEM[6991] <= 8'h62;
ROM_MEM[6992] <= 8'h80;
ROM_MEM[6993] <= 8'h62;
ROM_MEM[6994] <= 8'h80;
ROM_MEM[6995] <= 8'h62;
ROM_MEM[6996] <= 8'h90;
ROM_MEM[6997] <= 8'h62;
ROM_MEM[6998] <= 8'h90;
ROM_MEM[6999] <= 8'h62;
ROM_MEM[7000] <= 8'hA0;
ROM_MEM[7001] <= 8'h62;
ROM_MEM[7002] <= 8'hA0;
ROM_MEM[7003] <= 8'h67;
ROM_MEM[7004] <= 8'h80;
ROM_MEM[7005] <= 8'h62;
ROM_MEM[7006] <= 8'hA0;
ROM_MEM[7007] <= 8'h67;
ROM_MEM[7008] <= 8'h90;
ROM_MEM[7009] <= 8'h62;
ROM_MEM[7010] <= 8'hA0;
ROM_MEM[7011] <= 8'h67;
ROM_MEM[7012] <= 8'hA0;
ROM_MEM[7013] <= 8'h62;
ROM_MEM[7014] <= 8'hA0;
ROM_MEM[7015] <= 8'h67;
ROM_MEM[7016] <= 8'hC0;
ROM_MEM[7017] <= 8'h62;
ROM_MEM[7018] <= 8'hA0;
ROM_MEM[7019] <= 8'h66;
ROM_MEM[7020] <= 8'hA0;
ROM_MEM[7021] <= 8'h66;
ROM_MEM[7022] <= 8'hA0;
ROM_MEM[7023] <= 8'h66;
ROM_MEM[7024] <= 8'hA0;
ROM_MEM[7025] <= 8'h66;
ROM_MEM[7026] <= 8'hA0;
ROM_MEM[7027] <= 8'h66;
ROM_MEM[7028] <= 8'hA0;
ROM_MEM[7029] <= 8'h66;
ROM_MEM[7030] <= 8'hA0;
ROM_MEM[7031] <= 8'h66;
ROM_MEM[7032] <= 8'hA0;
ROM_MEM[7033] <= 8'h66;
ROM_MEM[7034] <= 8'hA0;
ROM_MEM[7035] <= 8'h86;
ROM_MEM[7036] <= 8'h01;
ROM_MEM[7037] <= 8'h97;
ROM_MEM[7038] <= 8'hA1;
ROM_MEM[7039] <= 8'hCC;
ROM_MEM[7040] <= 8'h00;
ROM_MEM[7041] <= 8'h01;
ROM_MEM[7042] <= 8'hDD;
ROM_MEM[7043] <= 8'h9F;
ROM_MEM[7044] <= 8'h39;
ROM_MEM[7045] <= 8'h96;
ROM_MEM[7046] <= 8'hA1;
ROM_MEM[7047] <= 8'h48;
ROM_MEM[7048] <= 8'h8E;
ROM_MEM[7049] <= 8'hBB;
ROM_MEM[7050] <= 8'h8E;
ROM_MEM[7051] <= 8'hAD;
ROM_MEM[7052] <= 8'h96;
ROM_MEM[7053] <= 8'h39;
ROM_MEM[7054] <= 8'hBB;
ROM_MEM[7055] <= 8'h8D;
ROM_MEM[7056] <= 8'hBB;
ROM_MEM[7057] <= 8'h98;
ROM_MEM[7058] <= 8'hBB;
ROM_MEM[7059] <= 8'hBB;
ROM_MEM[7060] <= 8'hBC;
ROM_MEM[7061] <= 8'h1E;
ROM_MEM[7062] <= 8'hBC;
ROM_MEM[7063] <= 8'h85;
ROM_MEM[7064] <= 8'hCC;
ROM_MEM[7065] <= 8'h64;
ROM_MEM[7066] <= 8'h80;
ROM_MEM[7067] <= 8'hCE;
ROM_MEM[7068] <= 8'h76;
ROM_MEM[7069] <= 8'hF0;
ROM_MEM[7070] <= 8'h9E;
ROM_MEM[7071] <= 8'h9F;
ROM_MEM[7072] <= 8'hBD;
ROM_MEM[7073] <= 8'hBC;
ROM_MEM[7074] <= 8'hAE;
ROM_MEM[7075] <= 8'hDC;
ROM_MEM[7076] <= 8'h9F;
ROM_MEM[7077] <= 8'hC3;
ROM_MEM[7078] <= 8'h00;
ROM_MEM[7079] <= 8'h02;
ROM_MEM[7080] <= 8'hDD;
ROM_MEM[7081] <= 8'h9F;
ROM_MEM[7082] <= 8'h10;
ROM_MEM[7083] <= 8'h83;
ROM_MEM[7084] <= 8'h00;
ROM_MEM[7085] <= 8'h3F;
ROM_MEM[7086] <= 8'h24;
ROM_MEM[7087] <= 8'h0A;
ROM_MEM[7088] <= 8'hCC;
ROM_MEM[7089] <= 8'h00;
ROM_MEM[7090] <= 8'h01;
ROM_MEM[7091] <= 8'hDD;
ROM_MEM[7092] <= 8'h9F;
ROM_MEM[7093] <= 8'h0C;
ROM_MEM[7094] <= 8'hA1;
ROM_MEM[7095] <= 8'hBD;
ROM_MEM[7096] <= 8'hBD;
ROM_MEM[7097] <= 8'hB7;
ROM_MEM[7098] <= 8'h39;
ROM_MEM[7099] <= 8'h9E;
ROM_MEM[7100] <= 8'h9F;
ROM_MEM[7101] <= 8'hCC;
ROM_MEM[7102] <= 8'h61;
ROM_MEM[7103] <= 8'hFF;
ROM_MEM[7104] <= 8'hCE;
ROM_MEM[7105] <= 8'h76;
ROM_MEM[7106] <= 8'hF0;
ROM_MEM[7107] <= 8'hBD;
ROM_MEM[7108] <= 8'hBC;
ROM_MEM[7109] <= 8'hAE;
ROM_MEM[7110] <= 8'hDC;
ROM_MEM[7111] <= 8'h9F;
ROM_MEM[7112] <= 8'hC3;
ROM_MEM[7113] <= 8'h00;
ROM_MEM[7114] <= 8'h02;
ROM_MEM[7115] <= 8'hDD;
ROM_MEM[7116] <= 8'h9F;
ROM_MEM[7117] <= 8'h10;
ROM_MEM[7118] <= 8'h83;
ROM_MEM[7119] <= 8'h00;
ROM_MEM[7120] <= 8'h3F;
ROM_MEM[7121] <= 8'h24;
ROM_MEM[7122] <= 8'h38;
ROM_MEM[7123] <= 8'hC6;
ROM_MEM[7124] <= 8'h3F;
ROM_MEM[7125] <= 8'hD0;
ROM_MEM[7126] <= 8'hA0;
ROM_MEM[7127] <= 8'h4F;
ROM_MEM[7128] <= 8'h1F;
ROM_MEM[7129] <= 8'h01;
ROM_MEM[7130] <= 8'hCC;
ROM_MEM[7131] <= 8'h64;
ROM_MEM[7132] <= 8'hFF;
ROM_MEM[7133] <= 8'hBD;
ROM_MEM[7134] <= 8'hBC;
ROM_MEM[7135] <= 8'hAE;
ROM_MEM[7136] <= 8'hDC;
ROM_MEM[7137] <= 8'h9F;
ROM_MEM[7138] <= 8'h58;
ROM_MEM[7139] <= 8'h49;
ROM_MEM[7140] <= 8'h58;
ROM_MEM[7141] <= 8'h49;
ROM_MEM[7142] <= 8'h58;
ROM_MEM[7143] <= 8'h49;
ROM_MEM[7144] <= 8'h43;
ROM_MEM[7145] <= 8'h53;
ROM_MEM[7146] <= 8'h2B;
ROM_MEM[7147] <= 8'h03;
ROM_MEM[7148] <= 8'h4A;
ROM_MEM[7149] <= 8'hCA;
ROM_MEM[7150] <= 8'h80;
ROM_MEM[7151] <= 8'hC3;
ROM_MEM[7152] <= 8'h76;
ROM_MEM[7153] <= 8'h70;
ROM_MEM[7154] <= 8'h5D;
ROM_MEM[7155] <= 8'h2B;
ROM_MEM[7156] <= 8'h03;
ROM_MEM[7157] <= 8'h4A;
ROM_MEM[7158] <= 8'hC4;
ROM_MEM[7159] <= 8'h7F;
ROM_MEM[7160] <= 8'h1F;
ROM_MEM[7161] <= 8'h03;
ROM_MEM[7162] <= 8'hDC;
ROM_MEM[7163] <= 8'h9F;
ROM_MEM[7164] <= 8'h54;
ROM_MEM[7165] <= 8'h54;
ROM_MEM[7166] <= 8'hC4;
ROM_MEM[7167] <= 8'h07;
ROM_MEM[7168] <= 8'hC8;
ROM_MEM[7169] <= 8'h07;
ROM_MEM[7170] <= 8'h5C;
ROM_MEM[7171] <= 8'h1F;
ROM_MEM[7172] <= 8'h01;
ROM_MEM[7173] <= 8'hCC;
ROM_MEM[7174] <= 8'h64;
ROM_MEM[7175] <= 8'hFF;
ROM_MEM[7176] <= 8'hBD;
ROM_MEM[7177] <= 8'hBC;
ROM_MEM[7178] <= 8'hC8;
ROM_MEM[7179] <= 8'hDC;
ROM_MEM[7180] <= 8'h9F;
ROM_MEM[7181] <= 8'h10;
ROM_MEM[7182] <= 8'h83;
ROM_MEM[7183] <= 8'h00;
ROM_MEM[7184] <= 8'h3F;
ROM_MEM[7185] <= 8'h25;
ROM_MEM[7186] <= 8'h0A;
ROM_MEM[7187] <= 8'hCC;
ROM_MEM[7188] <= 8'h00;
ROM_MEM[7189] <= 8'h01;
ROM_MEM[7190] <= 8'hDD;
ROM_MEM[7191] <= 8'h9F;
ROM_MEM[7192] <= 8'h0C;
ROM_MEM[7193] <= 8'hA1;
ROM_MEM[7194] <= 8'hBD;
ROM_MEM[7195] <= 8'hBD;
ROM_MEM[7196] <= 8'hB7;
ROM_MEM[7197] <= 8'h39;
ROM_MEM[7198] <= 8'h9E;
ROM_MEM[7199] <= 8'h9F;
ROM_MEM[7200] <= 8'hCC;
ROM_MEM[7201] <= 8'h67;
ROM_MEM[7202] <= 8'hFF;
ROM_MEM[7203] <= 8'hCE;
ROM_MEM[7204] <= 8'h76;
ROM_MEM[7205] <= 8'h70;
ROM_MEM[7206] <= 8'hBD;
ROM_MEM[7207] <= 8'hBC;
ROM_MEM[7208] <= 8'hAE;
ROM_MEM[7209] <= 8'hDC;
ROM_MEM[7210] <= 8'h9F;
ROM_MEM[7211] <= 8'hC3;
ROM_MEM[7212] <= 8'h00;
ROM_MEM[7213] <= 8'h03;
ROM_MEM[7214] <= 8'hDD;
ROM_MEM[7215] <= 8'h9F;
ROM_MEM[7216] <= 8'h10;
ROM_MEM[7217] <= 8'h83;
ROM_MEM[7218] <= 8'h00;
ROM_MEM[7219] <= 8'h3F;
ROM_MEM[7220] <= 8'h24;
ROM_MEM[7221] <= 8'h0D;
ROM_MEM[7222] <= 8'hC6;
ROM_MEM[7223] <= 8'h3F;
ROM_MEM[7224] <= 8'hD0;
ROM_MEM[7225] <= 8'hA0;
ROM_MEM[7226] <= 8'h4F;
ROM_MEM[7227] <= 8'h1F;
ROM_MEM[7228] <= 8'h01;
ROM_MEM[7229] <= 8'hCC;
ROM_MEM[7230] <= 8'h61;
ROM_MEM[7231] <= 8'hFF;
ROM_MEM[7232] <= 8'hBD;
ROM_MEM[7233] <= 8'hBC;
ROM_MEM[7234] <= 8'hAE;
ROM_MEM[7235] <= 8'hDC;
ROM_MEM[7236] <= 8'h9F;
ROM_MEM[7237] <= 8'h10;
ROM_MEM[7238] <= 8'h83;
ROM_MEM[7239] <= 8'h00;
ROM_MEM[7240] <= 8'h3F;
ROM_MEM[7241] <= 8'h24;
ROM_MEM[7242] <= 8'h27;
ROM_MEM[7243] <= 8'h58;
ROM_MEM[7244] <= 8'h49;
ROM_MEM[7245] <= 8'h58;
ROM_MEM[7246] <= 8'h49;
ROM_MEM[7247] <= 8'h58;
ROM_MEM[7248] <= 8'h49;
ROM_MEM[7249] <= 8'h43;
ROM_MEM[7250] <= 8'h53;
ROM_MEM[7251] <= 8'h2B;
ROM_MEM[7252] <= 8'h03;
ROM_MEM[7253] <= 8'h4A;
ROM_MEM[7254] <= 8'hCA;
ROM_MEM[7255] <= 8'h80;
ROM_MEM[7256] <= 8'hC3;
ROM_MEM[7257] <= 8'h76;
ROM_MEM[7258] <= 8'h70;
ROM_MEM[7259] <= 8'h5D;
ROM_MEM[7260] <= 8'h2B;
ROM_MEM[7261] <= 8'h03;
ROM_MEM[7262] <= 8'h4A;
ROM_MEM[7263] <= 8'hC4;
ROM_MEM[7264] <= 8'h7F;
ROM_MEM[7265] <= 8'h1F;
ROM_MEM[7266] <= 8'h03;
ROM_MEM[7267] <= 8'hDC;
ROM_MEM[7268] <= 8'h9F;
ROM_MEM[7269] <= 8'hC4;
ROM_MEM[7270] <= 8'h0F;
ROM_MEM[7271] <= 8'hC8;
ROM_MEM[7272] <= 8'h0F;
ROM_MEM[7273] <= 8'h5C;
ROM_MEM[7274] <= 8'h1F;
ROM_MEM[7275] <= 8'h01;
ROM_MEM[7276] <= 8'hCC;
ROM_MEM[7277] <= 8'h61;
ROM_MEM[7278] <= 8'hFF;
ROM_MEM[7279] <= 8'hBD;
ROM_MEM[7280] <= 8'hBC;
ROM_MEM[7281] <= 8'hC8;
ROM_MEM[7282] <= 8'hDC;
ROM_MEM[7283] <= 8'h9F;
ROM_MEM[7284] <= 8'h10;
ROM_MEM[7285] <= 8'h83;
ROM_MEM[7286] <= 8'h00;
ROM_MEM[7287] <= 8'h50;
ROM_MEM[7288] <= 8'h25;
ROM_MEM[7289] <= 8'h0A;
ROM_MEM[7290] <= 8'hCC;
ROM_MEM[7291] <= 8'h00;
ROM_MEM[7292] <= 8'h80;
ROM_MEM[7293] <= 8'hDD;
ROM_MEM[7294] <= 8'h9F;
ROM_MEM[7295] <= 8'h0C;
ROM_MEM[7296] <= 8'hA1;
ROM_MEM[7297] <= 8'hBD;
ROM_MEM[7298] <= 8'hBD;
ROM_MEM[7299] <= 8'hB7;
ROM_MEM[7300] <= 8'h39;
ROM_MEM[7301] <= 8'hDC;
ROM_MEM[7302] <= 8'h9F;
ROM_MEM[7303] <= 8'h83;
ROM_MEM[7304] <= 8'h00;
ROM_MEM[7305] <= 8'h04;
ROM_MEM[7306] <= 8'hDD;
ROM_MEM[7307] <= 8'h9F;
ROM_MEM[7308] <= 8'h10;
ROM_MEM[7309] <= 8'h83;
ROM_MEM[7310] <= 8'h00;
ROM_MEM[7311] <= 8'h08;
ROM_MEM[7312] <= 8'h25;
ROM_MEM[7313] <= 8'h17;
ROM_MEM[7314] <= 8'hC3;
ROM_MEM[7315] <= 8'h75;
ROM_MEM[7316] <= 8'h00;
ROM_MEM[7317] <= 8'h1F;
ROM_MEM[7318] <= 8'h03;
ROM_MEM[7319] <= 8'hDC;
ROM_MEM[7320] <= 8'h9F;
ROM_MEM[7321] <= 8'h44;
ROM_MEM[7322] <= 8'h56;
ROM_MEM[7323] <= 8'hC4;
ROM_MEM[7324] <= 8'h3F;
ROM_MEM[7325] <= 8'hC8;
ROM_MEM[7326] <= 8'h3F;
ROM_MEM[7327] <= 8'h1F;
ROM_MEM[7328] <= 8'h01;
ROM_MEM[7329] <= 8'hCC;
ROM_MEM[7330] <= 8'h67;
ROM_MEM[7331] <= 8'hFF;
ROM_MEM[7332] <= 8'hBD;
ROM_MEM[7333] <= 8'hBC;
ROM_MEM[7334] <= 8'hC8;
ROM_MEM[7335] <= 8'h20;
ROM_MEM[7336] <= 8'h04;
ROM_MEM[7337] <= 8'h86;
ROM_MEM[7338] <= 8'h00;
ROM_MEM[7339] <= 8'h97;
ROM_MEM[7340] <= 8'hA1;
ROM_MEM[7341] <= 8'h39;
ROM_MEM[7342] <= 8'hED;
ROM_MEM[7343] <= 8'hA1;
ROM_MEM[7344] <= 8'hCC;
ROM_MEM[7345] <= 8'h1F;
ROM_MEM[7346] <= 8'h98;
ROM_MEM[7347] <= 8'hED;
ROM_MEM[7348] <= 8'hA1;
ROM_MEM[7349] <= 8'hCC;
ROM_MEM[7350] <= 8'h00;
ROM_MEM[7351] <= 8'h00;
ROM_MEM[7352] <= 8'hED;
ROM_MEM[7353] <= 8'hA1;
ROM_MEM[7354] <= 8'hEF;
ROM_MEM[7355] <= 8'hA1;
ROM_MEM[7356] <= 8'hCC;
ROM_MEM[7357] <= 8'hBD;
ROM_MEM[7358] <= 8'h69;
ROM_MEM[7359] <= 8'hED;
ROM_MEM[7360] <= 8'hA1;
ROM_MEM[7361] <= 8'h33;
ROM_MEM[7362] <= 8'h5E;
ROM_MEM[7363] <= 8'h30;
ROM_MEM[7364] <= 8'h1F;
ROM_MEM[7365] <= 8'h26;
ROM_MEM[7366] <= 8'hE9;
ROM_MEM[7367] <= 8'h39;
ROM_MEM[7368] <= 8'hED;
ROM_MEM[7369] <= 8'hA1;
ROM_MEM[7370] <= 8'hCC;
ROM_MEM[7371] <= 8'h1F;
ROM_MEM[7372] <= 8'h98;
ROM_MEM[7373] <= 8'hED;
ROM_MEM[7374] <= 8'hA1;
ROM_MEM[7375] <= 8'hCC;
ROM_MEM[7376] <= 8'h00;
ROM_MEM[7377] <= 8'h00;
ROM_MEM[7378] <= 8'hED;
ROM_MEM[7379] <= 8'hA1;
ROM_MEM[7380] <= 8'hEF;
ROM_MEM[7381] <= 8'hA1;
ROM_MEM[7382] <= 8'hCC;
ROM_MEM[7383] <= 8'hBD;
ROM_MEM[7384] <= 8'h69;
ROM_MEM[7385] <= 8'hED;
ROM_MEM[7386] <= 8'hA1;
ROM_MEM[7387] <= 8'h1F;
ROM_MEM[7388] <= 8'h30;
ROM_MEM[7389] <= 8'h83;
ROM_MEM[7390] <= 8'h00;
ROM_MEM[7391] <= 8'h04;
ROM_MEM[7392] <= 8'hC4;
ROM_MEM[7393] <= 8'h7F;
ROM_MEM[7394] <= 8'h1F;
ROM_MEM[7395] <= 8'h03;
ROM_MEM[7396] <= 8'h30;
ROM_MEM[7397] <= 8'h1F;
ROM_MEM[7398] <= 8'h26;
ROM_MEM[7399] <= 8'hE2;
ROM_MEM[7400] <= 8'h39;
ROM_MEM[7401] <= 8'hC6;
ROM_MEM[7402] <= 8'h0E;
ROM_MEM[7403] <= 8'h7D;
ROM_MEM[7404] <= 8'h44;
ROM_MEM[7405] <= 8'h01;
ROM_MEM[7406] <= 8'h2A;
ROM_MEM[7407] <= 8'h05;
ROM_MEM[7408] <= 8'h5A;
ROM_MEM[7409] <= 8'h26;
ROM_MEM[7410] <= 8'hF8;
ROM_MEM[7411] <= 8'h86;
ROM_MEM[7412] <= 8'h00;
ROM_MEM[7413] <= 8'hB7;
ROM_MEM[7414] <= 8'h44;
ROM_MEM[7415] <= 8'h00;
ROM_MEM[7416] <= 8'h39;
ROM_MEM[7417] <= 8'h86;
ROM_MEM[7418] <= 8'h01;
ROM_MEM[7419] <= 8'h7E;
ROM_MEM[7420] <= 8'hBC;
ROM_MEM[7421] <= 8'hE9;
ROM_MEM[7422] <= 8'h86;
ROM_MEM[7423] <= 8'h02;
ROM_MEM[7424] <= 8'h7E;
ROM_MEM[7425] <= 8'hBC;
ROM_MEM[7426] <= 8'hE9;
ROM_MEM[7427] <= 8'h86;
ROM_MEM[7428] <= 8'h03;
ROM_MEM[7429] <= 8'h7E;
ROM_MEM[7430] <= 8'hBC;
ROM_MEM[7431] <= 8'hE9;
ROM_MEM[7432] <= 8'h86;
ROM_MEM[7433] <= 8'h04;
ROM_MEM[7434] <= 8'h7E;
ROM_MEM[7435] <= 8'hBC;
ROM_MEM[7436] <= 8'hE9;
ROM_MEM[7437] <= 8'h86;
ROM_MEM[7438] <= 8'h05;
ROM_MEM[7439] <= 8'h7E;
ROM_MEM[7440] <= 8'hBC;
ROM_MEM[7441] <= 8'hE9;
ROM_MEM[7442] <= 8'h86;
ROM_MEM[7443] <= 8'h06;
ROM_MEM[7444] <= 8'h7E;
ROM_MEM[7445] <= 8'hBC;
ROM_MEM[7446] <= 8'hE9;
ROM_MEM[7447] <= 8'h86;
ROM_MEM[7448] <= 8'h07;
ROM_MEM[7449] <= 8'h7E;
ROM_MEM[7450] <= 8'hBC;
ROM_MEM[7451] <= 8'hE9;
ROM_MEM[7452] <= 8'h86;
ROM_MEM[7453] <= 8'h08;
ROM_MEM[7454] <= 8'h7E;
ROM_MEM[7455] <= 8'hBC;
ROM_MEM[7456] <= 8'hE9;
ROM_MEM[7457] <= 8'h86;
ROM_MEM[7458] <= 8'h09;
ROM_MEM[7459] <= 8'h7E;
ROM_MEM[7460] <= 8'hBC;
ROM_MEM[7461] <= 8'hE9;
ROM_MEM[7462] <= 8'h86;
ROM_MEM[7463] <= 8'h0A;
ROM_MEM[7464] <= 8'h7E;
ROM_MEM[7465] <= 8'hBC;
ROM_MEM[7466] <= 8'hE9;
ROM_MEM[7467] <= 8'h86;
ROM_MEM[7468] <= 8'h0B;
ROM_MEM[7469] <= 8'h7E;
ROM_MEM[7470] <= 8'hBC;
ROM_MEM[7471] <= 8'hE9;
ROM_MEM[7472] <= 8'h86;
ROM_MEM[7473] <= 8'h0C;
ROM_MEM[7474] <= 8'h7E;
ROM_MEM[7475] <= 8'hBC;
ROM_MEM[7476] <= 8'hE9;
ROM_MEM[7477] <= 8'h86;
ROM_MEM[7478] <= 8'h0D;
ROM_MEM[7479] <= 8'h7E;
ROM_MEM[7480] <= 8'hBC;
ROM_MEM[7481] <= 8'hE9;
ROM_MEM[7482] <= 8'h86;
ROM_MEM[7483] <= 8'h0E;
ROM_MEM[7484] <= 8'h7E;
ROM_MEM[7485] <= 8'hBC;
ROM_MEM[7486] <= 8'hE9;
ROM_MEM[7487] <= 8'h86;
ROM_MEM[7488] <= 8'h0F;
ROM_MEM[7489] <= 8'h7E;
ROM_MEM[7490] <= 8'hBC;
ROM_MEM[7491] <= 8'hE9;
ROM_MEM[7492] <= 8'h86;
ROM_MEM[7493] <= 8'h10;
ROM_MEM[7494] <= 8'h7E;
ROM_MEM[7495] <= 8'hBC;
ROM_MEM[7496] <= 8'hE9;
ROM_MEM[7497] <= 8'h86;
ROM_MEM[7498] <= 8'h11;
ROM_MEM[7499] <= 8'h7E;
ROM_MEM[7500] <= 8'hBC;
ROM_MEM[7501] <= 8'hE9;
ROM_MEM[7502] <= 8'h86;
ROM_MEM[7503] <= 8'h12;
ROM_MEM[7504] <= 8'h7E;
ROM_MEM[7505] <= 8'hBC;
ROM_MEM[7506] <= 8'hE9;
ROM_MEM[7507] <= 8'h86;
ROM_MEM[7508] <= 8'h13;
ROM_MEM[7509] <= 8'h7E;
ROM_MEM[7510] <= 8'hBC;
ROM_MEM[7511] <= 8'hE9;
ROM_MEM[7512] <= 8'h86;
ROM_MEM[7513] <= 8'h14;
ROM_MEM[7514] <= 8'h7E;
ROM_MEM[7515] <= 8'hBC;
ROM_MEM[7516] <= 8'hE9;
ROM_MEM[7517] <= 8'h86;
ROM_MEM[7518] <= 8'h15;
ROM_MEM[7519] <= 8'h7E;
ROM_MEM[7520] <= 8'hBC;
ROM_MEM[7521] <= 8'hE9;
ROM_MEM[7522] <= 8'h86;
ROM_MEM[7523] <= 8'h16;
ROM_MEM[7524] <= 8'h7E;
ROM_MEM[7525] <= 8'hBC;
ROM_MEM[7526] <= 8'hE9;
ROM_MEM[7527] <= 8'h86;
ROM_MEM[7528] <= 8'h17;
ROM_MEM[7529] <= 8'h7E;
ROM_MEM[7530] <= 8'hBC;
ROM_MEM[7531] <= 8'hE9;
ROM_MEM[7532] <= 8'h86;
ROM_MEM[7533] <= 8'h18;
ROM_MEM[7534] <= 8'h7E;
ROM_MEM[7535] <= 8'hBC;
ROM_MEM[7536] <= 8'hE9;
ROM_MEM[7537] <= 8'h86;
ROM_MEM[7538] <= 8'h19;
ROM_MEM[7539] <= 8'h7E;
ROM_MEM[7540] <= 8'hBC;
ROM_MEM[7541] <= 8'hE9;
ROM_MEM[7542] <= 8'h86;
ROM_MEM[7543] <= 8'h1A;
ROM_MEM[7544] <= 8'h7E;
ROM_MEM[7545] <= 8'hBC;
ROM_MEM[7546] <= 8'hE9;
ROM_MEM[7547] <= 8'h86;
ROM_MEM[7548] <= 8'h1B;
ROM_MEM[7549] <= 8'h7E;
ROM_MEM[7550] <= 8'hBC;
ROM_MEM[7551] <= 8'hE9;
ROM_MEM[7552] <= 8'h86;
ROM_MEM[7553] <= 8'h1C;
ROM_MEM[7554] <= 8'h7E;
ROM_MEM[7555] <= 8'hBC;
ROM_MEM[7556] <= 8'hE9;
ROM_MEM[7557] <= 8'h86;
ROM_MEM[7558] <= 8'h1D;
ROM_MEM[7559] <= 8'h7E;
ROM_MEM[7560] <= 8'hBC;
ROM_MEM[7561] <= 8'hE9;
ROM_MEM[7562] <= 8'h86;
ROM_MEM[7563] <= 8'h1E;
ROM_MEM[7564] <= 8'h7E;
ROM_MEM[7565] <= 8'hBC;
ROM_MEM[7566] <= 8'hE9;
ROM_MEM[7567] <= 8'h86;
ROM_MEM[7568] <= 8'h1F;
ROM_MEM[7569] <= 8'h7E;
ROM_MEM[7570] <= 8'hBC;
ROM_MEM[7571] <= 8'hE9;
ROM_MEM[7572] <= 8'h86;
ROM_MEM[7573] <= 8'h20;
ROM_MEM[7574] <= 8'h7E;
ROM_MEM[7575] <= 8'hBC;
ROM_MEM[7576] <= 8'hE9;
ROM_MEM[7577] <= 8'h86;
ROM_MEM[7578] <= 8'h21;
ROM_MEM[7579] <= 8'h7E;
ROM_MEM[7580] <= 8'hBC;
ROM_MEM[7581] <= 8'hE9;
ROM_MEM[7582] <= 8'h86;
ROM_MEM[7583] <= 8'h22;
ROM_MEM[7584] <= 8'h7E;
ROM_MEM[7585] <= 8'hBC;
ROM_MEM[7586] <= 8'hE9;
ROM_MEM[7587] <= 8'h86;
ROM_MEM[7588] <= 8'h23;
ROM_MEM[7589] <= 8'h7E;
ROM_MEM[7590] <= 8'hBC;
ROM_MEM[7591] <= 8'hE9;
ROM_MEM[7592] <= 8'h86;
ROM_MEM[7593] <= 8'h24;
ROM_MEM[7594] <= 8'h7E;
ROM_MEM[7595] <= 8'hBC;
ROM_MEM[7596] <= 8'hE9;
ROM_MEM[7597] <= 8'h86;
ROM_MEM[7598] <= 8'h25;
ROM_MEM[7599] <= 8'h7E;
ROM_MEM[7600] <= 8'hBC;
ROM_MEM[7601] <= 8'hE9;
ROM_MEM[7602] <= 8'h86;
ROM_MEM[7603] <= 8'h26;
ROM_MEM[7604] <= 8'h7E;
ROM_MEM[7605] <= 8'hBC;
ROM_MEM[7606] <= 8'hE9;
ROM_MEM[7607] <= 8'h86;
ROM_MEM[7608] <= 8'h27;
ROM_MEM[7609] <= 8'h7E;
ROM_MEM[7610] <= 8'hBC;
ROM_MEM[7611] <= 8'hE9;
ROM_MEM[7612] <= 8'h86;
ROM_MEM[7613] <= 8'h28;
ROM_MEM[7614] <= 8'h7E;
ROM_MEM[7615] <= 8'hBC;
ROM_MEM[7616] <= 8'hE9;
ROM_MEM[7617] <= 8'h86;
ROM_MEM[7618] <= 8'h29;
ROM_MEM[7619] <= 8'h7E;
ROM_MEM[7620] <= 8'hBC;
ROM_MEM[7621] <= 8'hE9;
ROM_MEM[7622] <= 8'h86;
ROM_MEM[7623] <= 8'h2A;
ROM_MEM[7624] <= 8'h7E;
ROM_MEM[7625] <= 8'hBC;
ROM_MEM[7626] <= 8'hE9;
ROM_MEM[7627] <= 8'h86;
ROM_MEM[7628] <= 8'h2B;
ROM_MEM[7629] <= 8'h7E;
ROM_MEM[7630] <= 8'hBC;
ROM_MEM[7631] <= 8'hE9;
ROM_MEM[7632] <= 8'h86;
ROM_MEM[7633] <= 8'h2C;
ROM_MEM[7634] <= 8'h7E;
ROM_MEM[7635] <= 8'hBC;
ROM_MEM[7636] <= 8'hE9;
ROM_MEM[7637] <= 8'h86;
ROM_MEM[7638] <= 8'h2D;
ROM_MEM[7639] <= 8'h7E;
ROM_MEM[7640] <= 8'hBC;
ROM_MEM[7641] <= 8'hE9;
ROM_MEM[7642] <= 8'h86;
ROM_MEM[7643] <= 8'h2E;
ROM_MEM[7644] <= 8'h7E;
ROM_MEM[7645] <= 8'hBC;
ROM_MEM[7646] <= 8'hE9;
ROM_MEM[7647] <= 8'h86;
ROM_MEM[7648] <= 8'h2F;
ROM_MEM[7649] <= 8'h7E;
ROM_MEM[7650] <= 8'hBC;
ROM_MEM[7651] <= 8'hE9;
ROM_MEM[7652] <= 8'h86;
ROM_MEM[7653] <= 8'h30;
ROM_MEM[7654] <= 8'h7E;
ROM_MEM[7655] <= 8'hBC;
ROM_MEM[7656] <= 8'hE9;
ROM_MEM[7657] <= 8'h86;
ROM_MEM[7658] <= 8'h31;
ROM_MEM[7659] <= 8'h7E;
ROM_MEM[7660] <= 8'hBC;
ROM_MEM[7661] <= 8'hE9;
ROM_MEM[7662] <= 8'h86;
ROM_MEM[7663] <= 8'h32;
ROM_MEM[7664] <= 8'h7E;
ROM_MEM[7665] <= 8'hBC;
ROM_MEM[7666] <= 8'hE9;
ROM_MEM[7667] <= 8'h86;
ROM_MEM[7668] <= 8'h33;
ROM_MEM[7669] <= 8'h7E;
ROM_MEM[7670] <= 8'hBC;
ROM_MEM[7671] <= 8'hE9;
ROM_MEM[7672] <= 8'h86;
ROM_MEM[7673] <= 8'h34;
ROM_MEM[7674] <= 8'h7E;
ROM_MEM[7675] <= 8'hBC;
ROM_MEM[7676] <= 8'hE9;
ROM_MEM[7677] <= 8'h86;
ROM_MEM[7678] <= 8'h35;
ROM_MEM[7679] <= 8'h7E;
ROM_MEM[7680] <= 8'hBC;
ROM_MEM[7681] <= 8'hE9;
ROM_MEM[7682] <= 8'h86;
ROM_MEM[7683] <= 8'h36;
ROM_MEM[7684] <= 8'h7E;
ROM_MEM[7685] <= 8'hBC;
ROM_MEM[7686] <= 8'hE9;
ROM_MEM[7687] <= 8'h86;
ROM_MEM[7688] <= 8'h37;
ROM_MEM[7689] <= 8'h7E;
ROM_MEM[7690] <= 8'hBC;
ROM_MEM[7691] <= 8'hE9;
ROM_MEM[7692] <= 8'h86;
ROM_MEM[7693] <= 8'h38;
ROM_MEM[7694] <= 8'h7E;
ROM_MEM[7695] <= 8'hBC;
ROM_MEM[7696] <= 8'hE9;
ROM_MEM[7697] <= 8'h86;
ROM_MEM[7698] <= 8'h39;
ROM_MEM[7699] <= 8'h7E;
ROM_MEM[7700] <= 8'hBC;
ROM_MEM[7701] <= 8'hE9;
ROM_MEM[7702] <= 8'h86;
ROM_MEM[7703] <= 8'h3A;
ROM_MEM[7704] <= 8'h7E;
ROM_MEM[7705] <= 8'hBC;
ROM_MEM[7706] <= 8'hE9;
ROM_MEM[7707] <= 8'h86;
ROM_MEM[7708] <= 8'h3B;
ROM_MEM[7709] <= 8'h7E;
ROM_MEM[7710] <= 8'hBC;
ROM_MEM[7711] <= 8'hE9;
ROM_MEM[7712] <= 8'h86;
ROM_MEM[7713] <= 8'h59;
ROM_MEM[7714] <= 8'hBD;
ROM_MEM[7715] <= 8'hD8;
ROM_MEM[7716] <= 8'hDF;
ROM_MEM[7717] <= 8'h4C;
ROM_MEM[7718] <= 8'h81;
ROM_MEM[7719] <= 8'h65;
ROM_MEM[7720] <= 8'h25;
ROM_MEM[7721] <= 8'hF8;
ROM_MEM[7722] <= 8'h86;
ROM_MEM[7723] <= 8'hD3;
ROM_MEM[7724] <= 8'hBD;
ROM_MEM[7725] <= 8'hD8;
ROM_MEM[7726] <= 8'hDF;
ROM_MEM[7727] <= 8'hCC;
ROM_MEM[7728] <= 8'h64;
ROM_MEM[7729] <= 8'h80;
ROM_MEM[7730] <= 8'hED;
ROM_MEM[7731] <= 8'hA1;
ROM_MEM[7732] <= 8'h8E;
ROM_MEM[7733] <= 8'h45;
ROM_MEM[7734] <= 8'h3C;
ROM_MEM[7735] <= 8'hCE;
ROM_MEM[7736] <= 8'hC7;
ROM_MEM[7737] <= 8'hBB;
ROM_MEM[7738] <= 8'hEC;
ROM_MEM[7739] <= 8'hC1;
ROM_MEM[7740] <= 8'hED;
ROM_MEM[7741] <= 8'hA1;
ROM_MEM[7742] <= 8'hCC;
ROM_MEM[7743] <= 8'h00;
ROM_MEM[7744] <= 8'h30;
ROM_MEM[7745] <= 8'hED;
ROM_MEM[7746] <= 8'hA1;
ROM_MEM[7747] <= 8'hFF;
ROM_MEM[7748] <= 8'h4A;
ROM_MEM[7749] <= 8'hFA;
ROM_MEM[7750] <= 8'hC6;
ROM_MEM[7751] <= 8'h05;
ROM_MEM[7752] <= 8'hD7;
ROM_MEM[7753] <= 8'hAD;
ROM_MEM[7754] <= 8'hC6;
ROM_MEM[7755] <= 8'h05;
ROM_MEM[7756] <= 8'hA6;
ROM_MEM[7757] <= 8'h80;
ROM_MEM[7758] <= 8'hBD;
ROM_MEM[7759] <= 8'hE7;
ROM_MEM[7760] <= 8'hAD;
ROM_MEM[7761] <= 8'h5A;
ROM_MEM[7762] <= 8'h2A;
ROM_MEM[7763] <= 8'hF8;
ROM_MEM[7764] <= 8'hCC;
ROM_MEM[7765] <= 8'h80;
ROM_MEM[7766] <= 8'h40;
ROM_MEM[7767] <= 8'hED;
ROM_MEM[7768] <= 8'hA1;
ROM_MEM[7769] <= 8'hFE;
ROM_MEM[7770] <= 8'h4A;
ROM_MEM[7771] <= 8'hFA;
ROM_MEM[7772] <= 8'h8C;
ROM_MEM[7773] <= 8'h45;
ROM_MEM[7774] <= 8'h54;
ROM_MEM[7775] <= 8'h25;
ROM_MEM[7776] <= 8'hD9;
ROM_MEM[7777] <= 8'hFC;
ROM_MEM[7778] <= 8'hC7;
ROM_MEM[7779] <= 8'hC1;
ROM_MEM[7780] <= 8'hED;
ROM_MEM[7781] <= 8'hA1;
ROM_MEM[7782] <= 8'hCC;
ROM_MEM[7783] <= 8'h01;
ROM_MEM[7784] <= 8'h3C;
ROM_MEM[7785] <= 8'hED;
ROM_MEM[7786] <= 8'hA1;
ROM_MEM[7787] <= 8'h86;
ROM_MEM[7788] <= 8'h01;
ROM_MEM[7789] <= 8'h97;
ROM_MEM[7790] <= 8'hAD;
ROM_MEM[7791] <= 8'hB6;
ROM_MEM[7792] <= 8'h45;
ROM_MEM[7793] <= 8'h88;
ROM_MEM[7794] <= 8'hBD;
ROM_MEM[7795] <= 8'hE7;
ROM_MEM[7796] <= 8'hAD;
ROM_MEM[7797] <= 8'hB6;
ROM_MEM[7798] <= 8'h45;
ROM_MEM[7799] <= 8'h89;
ROM_MEM[7800] <= 8'hBD;
ROM_MEM[7801] <= 8'hE7;
ROM_MEM[7802] <= 8'hAD;
ROM_MEM[7803] <= 8'hCC;
ROM_MEM[7804] <= 8'h80;
ROM_MEM[7805] <= 8'h40;
ROM_MEM[7806] <= 8'hED;
ROM_MEM[7807] <= 8'hA1;
ROM_MEM[7808] <= 8'h8E;
ROM_MEM[7809] <= 8'h45;
ROM_MEM[7810] <= 8'h48;
ROM_MEM[7811] <= 8'hBD;
ROM_MEM[7812] <= 8'hC6;
ROM_MEM[7813] <= 8'hD4;
ROM_MEM[7814] <= 8'hCE;
ROM_MEM[7815] <= 8'h4A;
ROM_MEM[7816] <= 8'hFE;
ROM_MEM[7817] <= 8'h8E;
ROM_MEM[7818] <= 8'h45;
ROM_MEM[7819] <= 8'h42;
ROM_MEM[7820] <= 8'hBD;
ROM_MEM[7821] <= 8'hC6;
ROM_MEM[7822] <= 8'hD7;
ROM_MEM[7823] <= 8'hB6;
ROM_MEM[7824] <= 8'h4A;
ROM_MEM[7825] <= 8'hFC;
ROM_MEM[7826] <= 8'hBB;
ROM_MEM[7827] <= 8'h4B;
ROM_MEM[7828] <= 8'h00;
ROM_MEM[7829] <= 8'h19;
ROM_MEM[7830] <= 8'hB7;
ROM_MEM[7831] <= 8'h4A;
ROM_MEM[7832] <= 8'hFC;
ROM_MEM[7833] <= 8'hB6;
ROM_MEM[7834] <= 8'h4A;
ROM_MEM[7835] <= 8'hFB;
ROM_MEM[7836] <= 8'hB9;
ROM_MEM[7837] <= 8'h4A;
ROM_MEM[7838] <= 8'hFF;
ROM_MEM[7839] <= 8'h19;
ROM_MEM[7840] <= 8'hB7;
ROM_MEM[7841] <= 8'h4A;
ROM_MEM[7842] <= 8'hFB;
ROM_MEM[7843] <= 8'hB6;
ROM_MEM[7844] <= 8'h4A;
ROM_MEM[7845] <= 8'hFA;
ROM_MEM[7846] <= 8'hB9;
ROM_MEM[7847] <= 8'h4A;
ROM_MEM[7848] <= 8'hFE;
ROM_MEM[7849] <= 8'h19;
ROM_MEM[7850] <= 8'hB7;
ROM_MEM[7851] <= 8'h4A;
ROM_MEM[7852] <= 8'hFA;
ROM_MEM[7853] <= 8'hFC;
ROM_MEM[7854] <= 8'hC7;
ROM_MEM[7855] <= 8'hC3;
ROM_MEM[7856] <= 8'hED;
ROM_MEM[7857] <= 8'hA1;
ROM_MEM[7858] <= 8'hCC;
ROM_MEM[7859] <= 8'h00;
ROM_MEM[7860] <= 8'h30;
ROM_MEM[7861] <= 8'hED;
ROM_MEM[7862] <= 8'hA1;
ROM_MEM[7863] <= 8'hC6;
ROM_MEM[7864] <= 8'h05;
ROM_MEM[7865] <= 8'hD7;
ROM_MEM[7866] <= 8'hAD;
ROM_MEM[7867] <= 8'hB6;
ROM_MEM[7868] <= 8'h4A;
ROM_MEM[7869] <= 8'hFA;
ROM_MEM[7870] <= 8'hBD;
ROM_MEM[7871] <= 8'hE7;
ROM_MEM[7872] <= 8'h90;
ROM_MEM[7873] <= 8'hB6;
ROM_MEM[7874] <= 8'h4A;
ROM_MEM[7875] <= 8'hFB;
ROM_MEM[7876] <= 8'hBD;
ROM_MEM[7877] <= 8'hE7;
ROM_MEM[7878] <= 8'h90;
ROM_MEM[7879] <= 8'hB6;
ROM_MEM[7880] <= 8'h4A;
ROM_MEM[7881] <= 8'hFC;
ROM_MEM[7882] <= 8'hBD;
ROM_MEM[7883] <= 8'hE7;
ROM_MEM[7884] <= 8'h90;
ROM_MEM[7885] <= 8'hCC;
ROM_MEM[7886] <= 8'h80;
ROM_MEM[7887] <= 8'h40;
ROM_MEM[7888] <= 8'hED;
ROM_MEM[7889] <= 8'hA1;
ROM_MEM[7890] <= 8'h8E;
ROM_MEM[7891] <= 8'h45;
ROM_MEM[7892] <= 8'h54;
ROM_MEM[7893] <= 8'hBD;
ROM_MEM[7894] <= 8'hC6;
ROM_MEM[7895] <= 8'hD4;
ROM_MEM[7896] <= 8'hBD;
ROM_MEM[7897] <= 8'hC0;
ROM_MEM[7898] <= 8'h87;
ROM_MEM[7899] <= 8'hFC;
ROM_MEM[7900] <= 8'hC7;
ROM_MEM[7901] <= 8'hC9;
ROM_MEM[7902] <= 8'hED;
ROM_MEM[7903] <= 8'hA1;
ROM_MEM[7904] <= 8'hCC;
ROM_MEM[7905] <= 8'h00;
ROM_MEM[7906] <= 8'h30;
ROM_MEM[7907] <= 8'hED;
ROM_MEM[7908] <= 8'hA1;
ROM_MEM[7909] <= 8'hC6;
ROM_MEM[7910] <= 8'h07;
ROM_MEM[7911] <= 8'hD7;
ROM_MEM[7912] <= 8'hAD;
ROM_MEM[7913] <= 8'hB6;
ROM_MEM[7914] <= 8'h4A;
ROM_MEM[7915] <= 8'hFA;
ROM_MEM[7916] <= 8'hBD;
ROM_MEM[7917] <= 8'hE7;
ROM_MEM[7918] <= 8'h90;
ROM_MEM[7919] <= 8'hB6;
ROM_MEM[7920] <= 8'h4A;
ROM_MEM[7921] <= 8'hFB;
ROM_MEM[7922] <= 8'hBD;
ROM_MEM[7923] <= 8'hE7;
ROM_MEM[7924] <= 8'h90;
ROM_MEM[7925] <= 8'hB6;
ROM_MEM[7926] <= 8'h4A;
ROM_MEM[7927] <= 8'hFC;
ROM_MEM[7928] <= 8'hBD;
ROM_MEM[7929] <= 8'hE7;
ROM_MEM[7930] <= 8'h90;
ROM_MEM[7931] <= 8'hB6;
ROM_MEM[7932] <= 8'h4A;
ROM_MEM[7933] <= 8'hFD;
ROM_MEM[7934] <= 8'hBD;
ROM_MEM[7935] <= 8'hE7;
ROM_MEM[7936] <= 8'h90;
ROM_MEM[7937] <= 8'hCC;
ROM_MEM[7938] <= 8'h80;
ROM_MEM[7939] <= 8'h40;
ROM_MEM[7940] <= 8'hED;
ROM_MEM[7941] <= 8'hA1;
ROM_MEM[7942] <= 8'h8E;
ROM_MEM[7943] <= 8'h45;
ROM_MEM[7944] <= 8'h5C;
ROM_MEM[7945] <= 8'hBD;
ROM_MEM[7946] <= 8'hC6;
ROM_MEM[7947] <= 8'hD4;
ROM_MEM[7948] <= 8'hBD;
ROM_MEM[7949] <= 8'hC0;
ROM_MEM[7950] <= 8'h87;
ROM_MEM[7951] <= 8'hFC;
ROM_MEM[7952] <= 8'hC7;
ROM_MEM[7953] <= 8'hCB;
ROM_MEM[7954] <= 8'hED;
ROM_MEM[7955] <= 8'hA1;
ROM_MEM[7956] <= 8'hCC;
ROM_MEM[7957] <= 8'h00;
ROM_MEM[7958] <= 8'h30;
ROM_MEM[7959] <= 8'hED;
ROM_MEM[7960] <= 8'hA1;
ROM_MEM[7961] <= 8'hC6;
ROM_MEM[7962] <= 8'h07;
ROM_MEM[7963] <= 8'hD7;
ROM_MEM[7964] <= 8'hAD;
ROM_MEM[7965] <= 8'hB6;
ROM_MEM[7966] <= 8'h4A;
ROM_MEM[7967] <= 8'hFA;
ROM_MEM[7968] <= 8'hBD;
ROM_MEM[7969] <= 8'hE7;
ROM_MEM[7970] <= 8'h90;
ROM_MEM[7971] <= 8'hB6;
ROM_MEM[7972] <= 8'h4A;
ROM_MEM[7973] <= 8'hFB;
ROM_MEM[7974] <= 8'hBD;
ROM_MEM[7975] <= 8'hE7;
ROM_MEM[7976] <= 8'h90;
ROM_MEM[7977] <= 8'hB6;
ROM_MEM[7978] <= 8'h4A;
ROM_MEM[7979] <= 8'hFC;
ROM_MEM[7980] <= 8'hBD;
ROM_MEM[7981] <= 8'hE7;
ROM_MEM[7982] <= 8'h90;
ROM_MEM[7983] <= 8'hB6;
ROM_MEM[7984] <= 8'h4A;
ROM_MEM[7985] <= 8'hFD;
ROM_MEM[7986] <= 8'hBD;
ROM_MEM[7987] <= 8'hE7;
ROM_MEM[7988] <= 8'h90;
ROM_MEM[7989] <= 8'hCC;
ROM_MEM[7990] <= 8'h80;
ROM_MEM[7991] <= 8'h40;
ROM_MEM[7992] <= 8'hED;
ROM_MEM[7993] <= 8'hA1;
ROM_MEM[7994] <= 8'h8E;
ROM_MEM[7995] <= 8'h45;
ROM_MEM[7996] <= 8'h4C;
ROM_MEM[7997] <= 8'hBD;
ROM_MEM[7998] <= 8'hC6;
ROM_MEM[7999] <= 8'hD4;
ROM_MEM[8000] <= 8'h7F;
ROM_MEM[8001] <= 8'h4A;
ROM_MEM[8002] <= 8'hFA;
ROM_MEM[8003] <= 8'hB6;
ROM_MEM[8004] <= 8'h4A;
ROM_MEM[8005] <= 8'hFB;
ROM_MEM[8006] <= 8'hBA;
ROM_MEM[8007] <= 8'h4A;
ROM_MEM[8008] <= 8'hFC;
ROM_MEM[8009] <= 8'hBA;
ROM_MEM[8010] <= 8'h4A;
ROM_MEM[8011] <= 8'hFD;
ROM_MEM[8012] <= 8'h27;
ROM_MEM[8013] <= 8'h2E;
ROM_MEM[8014] <= 8'h8E;
ROM_MEM[8015] <= 8'h45;
ROM_MEM[8016] <= 8'h54;
ROM_MEM[8017] <= 8'hCE;
ROM_MEM[8018] <= 8'h4A;
ROM_MEM[8019] <= 8'hFE;
ROM_MEM[8020] <= 8'hBD;
ROM_MEM[8021] <= 8'hC6;
ROM_MEM[8022] <= 8'hD7;
ROM_MEM[8023] <= 8'hBD;
ROM_MEM[8024] <= 8'hC0;
ROM_MEM[8025] <= 8'h2F;
ROM_MEM[8026] <= 8'hB6;
ROM_MEM[8027] <= 8'h4A;
ROM_MEM[8028] <= 8'hFA;
ROM_MEM[8029] <= 8'h84;
ROM_MEM[8030] <= 8'h0F;
ROM_MEM[8031] <= 8'h81;
ROM_MEM[8032] <= 8'h0F;
ROM_MEM[8033] <= 8'hB6;
ROM_MEM[8034] <= 8'h4A;
ROM_MEM[8035] <= 8'hFA;
ROM_MEM[8036] <= 8'h25;
ROM_MEM[8037] <= 8'h03;
ROM_MEM[8038] <= 8'h7C;
ROM_MEM[8039] <= 8'h4A;
ROM_MEM[8040] <= 8'hFA;
ROM_MEM[8041] <= 8'h44;
ROM_MEM[8042] <= 8'h44;
ROM_MEM[8043] <= 8'h44;
ROM_MEM[8044] <= 8'h44;
ROM_MEM[8045] <= 8'hBB;
ROM_MEM[8046] <= 8'h4A;
ROM_MEM[8047] <= 8'hFA;
ROM_MEM[8048] <= 8'hB7;
ROM_MEM[8049] <= 8'h4A;
ROM_MEM[8050] <= 8'hFA;
ROM_MEM[8051] <= 8'h84;
ROM_MEM[8052] <= 8'h0F;
ROM_MEM[8053] <= 8'h81;
ROM_MEM[8054] <= 8'h0F;
ROM_MEM[8055] <= 8'h25;
ROM_MEM[8056] <= 8'h03;
ROM_MEM[8057] <= 8'h7C;
ROM_MEM[8058] <= 8'h4A;
ROM_MEM[8059] <= 8'hFA;
ROM_MEM[8060] <= 8'hFC;
ROM_MEM[8061] <= 8'hC7;
ROM_MEM[8062] <= 8'hC5;
ROM_MEM[8063] <= 8'hED;
ROM_MEM[8064] <= 8'hA1;
ROM_MEM[8065] <= 8'hCC;
ROM_MEM[8066] <= 8'h00;
ROM_MEM[8067] <= 8'h30;
ROM_MEM[8068] <= 8'hED;
ROM_MEM[8069] <= 8'hA1;
ROM_MEM[8070] <= 8'hB6;
ROM_MEM[8071] <= 8'h4A;
ROM_MEM[8072] <= 8'hFA;
ROM_MEM[8073] <= 8'hBD;
ROM_MEM[8074] <= 8'hC7;
ROM_MEM[8075] <= 8'h0E;
ROM_MEM[8076] <= 8'hCC;
ROM_MEM[8077] <= 8'h80;
ROM_MEM[8078] <= 8'h40;
ROM_MEM[8079] <= 8'hED;
ROM_MEM[8080] <= 8'hA1;
ROM_MEM[8081] <= 8'h8E;
ROM_MEM[8082] <= 8'h45;
ROM_MEM[8083] <= 8'h5C;
ROM_MEM[8084] <= 8'hBD;
ROM_MEM[8085] <= 8'hC6;
ROM_MEM[8086] <= 8'hD4;
ROM_MEM[8087] <= 8'hB6;
ROM_MEM[8088] <= 8'h4A;
ROM_MEM[8089] <= 8'hFA;
ROM_MEM[8090] <= 8'hBA;
ROM_MEM[8091] <= 8'h4A;
ROM_MEM[8092] <= 8'hFB;
ROM_MEM[8093] <= 8'hBA;
ROM_MEM[8094] <= 8'h4A;
ROM_MEM[8095] <= 8'hFC;
ROM_MEM[8096] <= 8'hBA;
ROM_MEM[8097] <= 8'h4A;
ROM_MEM[8098] <= 8'hFD;
ROM_MEM[8099] <= 8'h27;
ROM_MEM[8100] <= 8'h0F;
ROM_MEM[8101] <= 8'h8E;
ROM_MEM[8102] <= 8'h45;
ROM_MEM[8103] <= 8'h56;
ROM_MEM[8104] <= 8'hCE;
ROM_MEM[8105] <= 8'h4A;
ROM_MEM[8106] <= 8'hFE;
ROM_MEM[8107] <= 8'hBD;
ROM_MEM[8108] <= 8'hC6;
ROM_MEM[8109] <= 8'hD7;
ROM_MEM[8110] <= 8'h7F;
ROM_MEM[8111] <= 8'h4B;
ROM_MEM[8112] <= 8'h01;
ROM_MEM[8113] <= 8'hBD;
ROM_MEM[8114] <= 8'hC0;
ROM_MEM[8115] <= 8'h2F;
ROM_MEM[8116] <= 8'hFC;
ROM_MEM[8117] <= 8'hC7;
ROM_MEM[8118] <= 8'hC7;
ROM_MEM[8119] <= 8'hED;
ROM_MEM[8120] <= 8'hA1;
ROM_MEM[8121] <= 8'hCC;
ROM_MEM[8122] <= 8'h00;
ROM_MEM[8123] <= 8'h30;
ROM_MEM[8124] <= 8'hED;
ROM_MEM[8125] <= 8'hA1;
ROM_MEM[8126] <= 8'h4F;
ROM_MEM[8127] <= 8'hF6;
ROM_MEM[8128] <= 8'h4A;
ROM_MEM[8129] <= 8'hFA;
ROM_MEM[8130] <= 8'h8E;
ROM_MEM[8131] <= 8'h00;
ROM_MEM[8132] <= 8'h10;
ROM_MEM[8133] <= 8'hBD;
ROM_MEM[8134] <= 8'h77;
ROM_MEM[8135] <= 8'h20;
ROM_MEM[8136] <= 8'hC6;
ROM_MEM[8137] <= 8'h01;
ROM_MEM[8138] <= 8'hD7;
ROM_MEM[8139] <= 8'hAD;
ROM_MEM[8140] <= 8'hB6;
ROM_MEM[8141] <= 8'h4A;
ROM_MEM[8142] <= 8'hD6;
ROM_MEM[8143] <= 8'hBD;
ROM_MEM[8144] <= 8'hE7;
ROM_MEM[8145] <= 8'h90;
ROM_MEM[8146] <= 8'hCC;
ROM_MEM[8147] <= 8'h80;
ROM_MEM[8148] <= 8'h40;
ROM_MEM[8149] <= 8'hED;
ROM_MEM[8150] <= 8'hA1;
ROM_MEM[8151] <= 8'hC6;
ROM_MEM[8152] <= 8'h11;
ROM_MEM[8153] <= 8'hF7;
ROM_MEM[8154] <= 8'h4A;
ROM_MEM[8155] <= 8'hFA;
ROM_MEM[8156] <= 8'hCE;
ROM_MEM[8157] <= 8'hC7;
ROM_MEM[8158] <= 8'hCD;
ROM_MEM[8159] <= 8'hFF;
ROM_MEM[8160] <= 8'h4A;
ROM_MEM[8161] <= 8'hFC;
ROM_MEM[8162] <= 8'hFE;
ROM_MEM[8163] <= 8'h4A;
ROM_MEM[8164] <= 8'hFC;
ROM_MEM[8165] <= 8'hEC;
ROM_MEM[8166] <= 8'hC1;
ROM_MEM[8167] <= 8'hED;
ROM_MEM[8168] <= 8'hA1;
ROM_MEM[8169] <= 8'h11;
ROM_MEM[8170] <= 8'h83;
ROM_MEM[8171] <= 8'hC7;
ROM_MEM[8172] <= 8'hE1;
ROM_MEM[8173] <= 8'h25;
ROM_MEM[8174] <= 8'h05;
ROM_MEM[8175] <= 8'hCC;
ROM_MEM[8176] <= 8'h1E;
ROM_MEM[8177] <= 8'hD4;
ROM_MEM[8178] <= 8'h20;
ROM_MEM[8179] <= 8'h03;
ROM_MEM[8180] <= 8'hCC;
ROM_MEM[8181] <= 8'h00;
ROM_MEM[8182] <= 8'h64;
ROM_MEM[8183] <= 8'hED;
ROM_MEM[8184] <= 8'hA1;
ROM_MEM[8185] <= 8'hFF;
ROM_MEM[8186] <= 8'h4A;
ROM_MEM[8187] <= 8'hFC;
ROM_MEM[8188] <= 8'h8E;
ROM_MEM[8189] <= 8'hC7;
ROM_MEM[8190] <= 8'hA3;
ROM_MEM[8191] <= 8'hF6;
    end
    
    reg [31:0] mem_reg;
    always @(posedge clk) begin
        data <= ROM_MEM[address];
    end
    
	
    
    
endmodule
