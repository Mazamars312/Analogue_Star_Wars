`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.05.2023 08:33:12
// Design Name: 
// Module Name: Vector_board
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module Vector_board(
//   input               	clk_12,
//   input               	clk_3,
//	input 					clk_1_5,
//	input 					clk_mpu,
//   input               	reset_n,
//    
//   input [15:0]        	main_cpu_address,
//   input [7:0]         	main_cpu_data_out,
//   input               	main_cpu_RnW,
//	 
//	input [23:0]			mpu_address,
//	input 					mpu_write,
//	input [3:0]				mpu_mask,
//	input 					mpu_request,
//	output reg  [31:0]	mpu_data_in,
//	input [31:0]			mpu_data_out,
//	output reg 				mpu_valid,
//    
//   output [7:0]        	V_data_out,
//   output reg          	VGHALT = 'b1,
//   input               	EVGRES_WR,
//   input               	EVGGO_WR
//   );
//    
    
//	wire [7:0]  cpu_vram_data_out;
//	wire [7:0]  cpu_vrom_data_out;
//
//	wire [31:0]  mpu_vram_data_out;
//	wire [31:0]  mpu_vrom_data_out;
//	
//	// MPS System
//	
//	reg EVGRES_WR_REG, EVGGO_WR_REG, mpu_request_reg;
//	
//	reg address_00;
//	reg address_01;
//	reg address_02;
//	reg address_03;
//	
////	wire mpu_write_VRAM = |{address_00, address_01, address_02} && mpu_write && mpu_request;
////	wire mpu_write_VROM =   address_03 && mpu_write && mpu_request_reg;
//	reg mpu_write_VRAM;
//	reg mpu_write_VROM;
//	always @(posedge clk_mpu) begin
//		address_00 <= (mpu_address[23:12] == 12'h000);
//		address_01 <= (mpu_address[23:12] == 12'h001);
//		address_02 <= (mpu_address[23:12] == 12'h002);
//		address_03 <= (mpu_address[23:12] == 12'h003);
//		mpu_write_VRAM <= |{address_00, address_01, address_02} && mpu_write && mpu_request_reg;
//		mpu_write_VROM <=   address_03 && mpu_write && mpu_request_reg;
//		mpu_request_reg <= mpu_request;
//	end
//	
//	
//
//	
//	wire EVGGO_WR_wire;
//	wire EVGRES_WR_wire;
//	
//	synch_3 s02(EVGGO_WR, EVGGO_WR_wire, clk_mpu);
//	synch_3 s03(EVGRES_WR, EVGRES_WR_wire, clk_mpu);
//	
//	always @(posedge clk_mpu or negedge reset_n) begin
//		if (~reset_n) begin
//			EVGRES_WR_REG	<=0; 
//			EVGGO_WR_REG	<=0;
//			VGHALT			<=0;
//		end
//		else begin
//		
//			EVGRES_WR_REG	<= EVGRES_WR_wire; 
//			EVGGO_WR_REG	<= EVGGO_WR_wire;
//			if (mpu_address[23:0] == 24'h00_4000 && mpu_request_reg && mpu_request) VGHALT <= mpu_data_out[0];
//			else begin
//				if (EVGRES_WR_wire && ~EVGRES_WR_REG) begin
//					VGHALT	<= 1;
//				end
//				if (EVGGO_WR_wire && ~EVGGO_WR_REG) begin
//					VGHALT	<= 0;
//				end
//			end
//		
//		end
//	end
	 
	 
    
//	assign V_data_out = main_cpu_address[13:12] == 'b11 ? cpu_vrom_data_out : cpu_vram_data_out;
//
//	wire vram_write = main_cpu_RnW && |{main_cpu_address[15:12] == 'b0000, main_cpu_address[15:12] == 'b0001, main_cpu_address[15:12] == 'b0010};
   // the sram port will be used for the Video buffer access and the System ROM/RAM access
	
	// 24'h01_0000			PROM 0 (16K)			0x4000	R/W
	// 24'h01_4000			PROM 1 (8K)				0x2000	R/W
	// 24'h01_6000			PROM 2 (8K)				0x2000	R/W
	// 24'h01_8000			PROM 3 (8K)				0x2000	R/W
	// 24'h01_A000			PROM 4 (8K)				0x2000	R/W
	// 24'h02_C000			Sound Rom 0 (8K)		0x2000	R/W
	// 24'h02_E000			Sound Rom 1 (8K)		0x2000	R/W
	// 24'h01_0000			matrix Rom 0 (1K)		0x400		R/W
	// 24'h01_0400			matrix Rom 1 (1K)		0x400		R/W
	// 24'h01_0800			matrix Rom 2 (1K)		0x400		R/W
	// 24'h01_0C00			matrix Rom 3 (1K)		0x400		R/W
	// 24'h00_0000			Vector Ram 0 (16K)	0x3000	R/W
	// 24'h00_3000			Vector Rom 0 (4K)		0x1000	R/W
	// 24'h00_4000			Vector_reg				0x4	R/W
	
	 
//	VRAM VRAM(
//	.clk_a		(clk_12),
//	.address_a	(main_cpu_address[13:0]),
//	.write_a		(vram_write),
//	.data_a		(main_cpu_data_out),
//	.q_a			(cpu_vram_data_out),
//
//	.clk_b		(clk_mpu),
//	.address_b	(mpu_address[13:2]),
//	.write_b		(mpu_write_VRAM),
//	.mask_b		(mpu_mask),
//	.data_b		({mpu_data_out[7:0], mpu_data_out[15:8], mpu_data_out[23:16],mpu_data_out[31:24]}),
//	.q_b			(mpu_vram_data_out),
//
//	);
// 
// 
//	VROM VROM(
//	.clk_a		(clk_12),
//	.address_a	(main_cpu_address[11:0]),
//	.q_a			(cpu_vrom_data_out),
//
//	.clk_b		(clk_mpu),
//	.address_b	(mpu_address[11:2]),
//	.write_b		(1'b0),
//	.mask_b		(mpu_mask),
//	.data_b		({mpu_data_out[7:0], mpu_data_out[15:8], mpu_data_out[23:16],mpu_data_out[31:24]}),
//	.q_b			(mpu_vrom_data_out),
//	);
 

    
//endmodule

module VRAM(
    input               clk_a,
    input      [13:0]  	address_a,
    input  		    		write_a,
    input  		[7:0]   	data_a,
    output reg [7:0]   	q_a,
	 
	 input               clk_b,
    input      [11:0]  	address_b,
    input  		    		write_b,
	 input		[3:0]		mask_b,
    input  		[31:0]   data_b,
    output 		[31:0]   q_b
    );
    
	 wire [31:0] q_a_reg;
	 reg [3:0] byteena_a;
	 
	 Vector_ram Vector_ram(
	.clock_a		(clk_a),
	.address_a	(address_a[13:2]),
	.wren_a		(write_a),
	.byteena_a	(byteena_a),
	.data_a		({4{data_a}}),
	.q_a			(q_a_reg),
	
	.clock_b		(clk_b),
	.wren_b		(write_b),
	.address_b	(address_b),
	.data_b		(data_b),
	.q_b			(q_b)
	);
	
	always @* begin
		case (address_a[1:0]) 
			2'b00 : q_a <= q_a_reg[31:24];
			2'b01 : q_a <= q_a_reg[23:16];
			2'b10 : q_a <= q_a_reg[15:8];
			2'b11 : q_a <= q_a_reg[7:0];
		endcase
	end
	
	always @* begin
		case (address_a[1:0]) 
			2'b00 	: byteena_a <= 4'b1000;
			2'b01 	: byteena_a <= 4'b0100;
			2'b10 	: byteena_a <= 4'b0010;
			default 	: byteena_a <= 4'b0001;
		endcase
	end
    
endmodule

module VROM(
    input               clk_a,
    input       [11:0]  address_a,
    output reg  [7:0]   q_a,
	 
	 
	 input               clk_b,
    input      [9:0]  	address_b,
    input  		    		write_b,
	 input		[3:0]		mask_b,
    input  		[31:0]   data_b,
    output reg [31:0]   q_b
    );
    
 reg [31:0] CPU_ROM_MEM [1023:0];
initial begin
CPU_ROM_MEM[0   ] <= 32'h1EECB87D;
CPU_ROM_MEM[1   ] <= 32'hB879B8B3;
CPU_ROM_MEM[2   ] <= 32'hB8B9B8BD;
CPU_ROM_MEM[3   ] <= 32'hB8C5B88F;
CPU_ROM_MEM[4   ] <= 32'hB8CAB8CF;
CPU_ROM_MEM[5   ] <= 32'hB8D4B8D7;
CPU_ROM_MEM[6   ] <= 32'hB82FB837;
CPU_ROM_MEM[7   ] <= 32'hB841B845;
CPU_ROM_MEM[8   ] <= 32'hB84CB84E;
CPU_ROM_MEM[9   ] <= 32'hB855B85A;
CPU_ROM_MEM[10  ] <= 32'hB85FB864;
CPU_ROM_MEM[11  ] <= 32'hB868B86E;
CPU_ROM_MEM[12  ] <= 32'hB872B876;
CPU_ROM_MEM[13  ] <= 32'hB879B87F;
CPU_ROM_MEM[14  ] <= 32'hB883B88B;
CPU_ROM_MEM[15  ] <= 32'hB88FB894;
CPU_ROM_MEM[16  ] <= 32'hB896B89C;
CPU_ROM_MEM[17  ] <= 32'hB8A0B8A5;
CPU_ROM_MEM[18  ] <= 32'hB8A9B8AF;
CPU_ROM_MEM[19  ] <= 32'hB8E6B8EA;
CPU_ROM_MEM[20  ] <= 32'hB8DCB8DF;
CPU_ROM_MEM[21  ] <= 32'hB870B8F3;
CPU_ROM_MEM[22  ] <= 32'hB8FFB90F;
CPU_ROM_MEM[23  ] <= 32'hC00048E0;
CPU_ROM_MEM[24  ] <= 32'h44E45CE4;
CPU_ROM_MEM[25  ] <= 32'h58E04518;
CPU_ROM_MEM[26  ] <= 32'h40E85B04;
CPU_ROM_MEM[27  ] <= 32'hC0004CE0;
CPU_ROM_MEM[28  ] <= 32'h40E55DE2;
CPU_ROM_MEM[29  ] <= 32'h5DFE40FB;
CPU_ROM_MEM[30  ] <= 32'h40065DE2;
CPU_ROM_MEM[31  ] <= 32'h5DFE40FA;
CPU_ROM_MEM[32  ] <= 32'hF87D4CE0;
CPU_ROM_MEM[33  ] <= 32'h40E85418;
CPU_ROM_MEM[34  ] <= 32'hF87040E5;
CPU_ROM_MEM[35  ] <= 32'h44E344E0;
CPU_ROM_MEM[36  ] <= 32'h44FD40FB;
CPU_ROM_MEM[37  ] <= 32'h54E0F87D;
CPU_ROM_MEM[38  ] <= 32'h40E84018;
CPU_ROM_MEM[39  ] <= 32'h460040E6;
CPU_ROM_MEM[40  ] <= 32'h5A1A4CE0;
CPU_ROM_MEM[41  ] <= 32'h40E8F89A;
CPU_ROM_MEM[42  ] <= 32'hC0004504;
CPU_ROM_MEM[43  ] <= 32'h40E45BE0;
CPU_ROM_MEM[44  ] <= 32'h4018F841;
CPU_ROM_MEM[45  ] <= 32'h4CE05A00;
CPU_ROM_MEM[46  ] <= 32'h40E85A00;
CPU_ROM_MEM[47  ] <= 32'hF89940E8;
CPU_ROM_MEM[48  ] <= 32'h4C1840E8;
CPU_ROM_MEM[49  ] <= 32'h401CF8B6;
CPU_ROM_MEM[50  ] <= 32'h44005CE4;
CPU_ROM_MEM[51  ] <= 32'h40E4F899;
CPU_ROM_MEM[52  ] <= 32'h4CE05A00;
CPU_ROM_MEM[53  ] <= 32'h46E85A18;
CPU_ROM_MEM[54  ] <= 32'h5AE8F8D2;
CPU_ROM_MEM[55  ] <= 32'h4C0054E0;
CPU_ROM_MEM[56  ] <= 32'h40E8F8D2;
CPU_ROM_MEM[57  ] <= 32'h4CE05CE4;
CPU_ROM_MEM[58  ] <= 32'h44E4F8D1;
CPU_ROM_MEM[59  ] <= 32'h4CE054E8;
CPU_ROM_MEM[60  ] <= 32'hF89940E8;
CPU_ROM_MEM[61  ] <= 32'h4CE05418;
CPU_ROM_MEM[62  ] <= 32'hF851400C;
CPU_ROM_MEM[63  ] <= 32'hC0004600;
CPU_ROM_MEM[64  ] <= 32'h40E846E0;
CPU_ROM_MEM[65  ] <= 32'hF87B4404;
CPU_ROM_MEM[66  ] <= 32'h5CE44018;
CPU_ROM_MEM[67  ] <= 32'h40E444E4;
CPU_ROM_MEM[68  ] <= 32'h48E05418;
CPU_ROM_MEM[69  ] <= 32'hF8514600;
CPU_ROM_MEM[70  ] <= 32'h5AE84018;
CPU_ROM_MEM[71  ] <= 32'hF87F4008;
CPU_ROM_MEM[72  ] <= 32'h46E04018;
CPU_ROM_MEM[73  ] <= 32'h46E0F8C0;
CPU_ROM_MEM[74  ] <= 32'h4C00F861;
CPU_ROM_MEM[75  ] <= 32'h4C0054E0;
CPU_ROM_MEM[76  ] <= 32'h40E84CE0;
CPU_ROM_MEM[77  ] <= 32'h5404C000;
CPU_ROM_MEM[78  ] <= 32'h4C0054E4;
CPU_ROM_MEM[79  ] <= 32'h4CE4F89A;
CPU_ROM_MEM[80  ] <= 32'h4C0054E0;
CPU_ROM_MEM[81  ] <= 32'h44E45CE4;
CPU_ROM_MEM[82  ] <= 32'hF8994CE8;
CPU_ROM_MEM[83  ] <= 32'h401854E8;
CPU_ROM_MEM[84  ] <= 32'hF8D24004;
CPU_ROM_MEM[85  ] <= 32'h48E044FC;
CPU_ROM_MEM[86  ] <= 32'h5C0444E4;
CPU_ROM_MEM[87  ] <= 32'hF89A4C00;
CPU_ROM_MEM[88  ] <= 32'h40E854F8;
CPU_ROM_MEM[89  ] <= 32'hF87040E8;
CPU_ROM_MEM[90  ] <= 32'h4A1A42E2;
CPU_ROM_MEM[91  ] <= 32'h54E04008;
CPU_ROM_MEM[92  ] <= 32'hC00046E0;
CPU_ROM_MEM[93  ] <= 32'h400846E0;
CPU_ROM_MEM[94  ] <= 32'hF8BF4008;
CPU_ROM_MEM[95  ] <= 32'h4CE04018;
CPU_ROM_MEM[96  ] <= 32'h40E85A18;
CPU_ROM_MEM[97  ] <= 32'h40E85A18;
CPU_ROM_MEM[98  ] <= 32'hF8704C00;
CPU_ROM_MEM[99  ] <= 32'h5AE040E8;
CPU_ROM_MEM[100 ] <= 32'h4600F8D1;
CPU_ROM_MEM[101 ] <= 32'h460040E8;
CPU_ROM_MEM[102 ] <= 32'h5AE04018;
CPU_ROM_MEM[103 ] <= 32'hF86E4C00;
CPU_ROM_MEM[104 ] <= 32'h40E854E0;
CPU_ROM_MEM[105 ] <= 32'h4004C000;
CPU_ROM_MEM[106 ] <= 32'h4CE05408;
CPU_ROM_MEM[107 ] <= 32'hF8BE4C00;
CPU_ROM_MEM[108 ] <= 32'h5AE040E8;
CPU_ROM_MEM[109 ] <= 32'h4618F8D0;
CPU_ROM_MEM[110 ] <= 32'h0000E000;
CPU_ROM_MEM[111 ] <= 32'hF87D4504;
CPU_ROM_MEM[112 ] <= 32'h0000E000;
CPU_ROM_MEM[113 ] <= 32'h5B000000;
CPU_ROM_MEM[114 ] <= 32'hE000F8B7;
CPU_ROM_MEM[115 ] <= 32'h4C05B8EE;
CPU_ROM_MEM[116 ] <= 32'h5407C000;
CPU_ROM_MEM[117 ] <= 32'h4002B8EE;
CPU_ROM_MEM[118 ] <= 32'h400AC000;
CPU_ROM_MEM[119 ] <= 32'h5BFE45E3;
CPU_ROM_MEM[120 ] <= 32'h0000FFFE;
CPU_ROM_MEM[121 ] <= 32'hC0004802;
CPU_ROM_MEM[122 ] <= 32'h44E0541E;
CPU_ROM_MEM[123 ] <= 32'h4CE65A1E;
CPU_ROM_MEM[124 ] <= 32'h40E45DE0;
CPU_ROM_MEM[125 ] <= 32'h40FB5DE0;
CPU_ROM_MEM[126 ] <= 32'h40E54004;
CPU_ROM_MEM[127 ] <= 32'hC0005D04;
CPU_ROM_MEM[128 ] <= 32'h45FC48E0;
CPU_ROM_MEM[129 ] <= 32'h45E440E8;
CPU_ROM_MEM[130 ] <= 32'h5B1F40FB;
CPU_ROM_MEM[131 ] <= 32'h57E040E5;
CPU_ROM_MEM[132 ] <= 32'h5C1940E8;
CPU_ROM_MEM[133 ] <= 32'h45E448E0;
CPU_ROM_MEM[134 ] <= 32'h45FC5100;
CPU_ROM_MEM[135 ] <= 32'hC0004601;
CPU_ROM_MEM[136 ] <= 32'h40E65A05;
CPU_ROM_MEM[137 ] <= 32'hC0005D1E;
CPU_ROM_MEM[138 ] <= 32'h45E15E03;
CPU_ROM_MEM[139 ] <= 32'hC00063FF;
CPU_ROM_MEM[140 ] <= 32'hC00061FF;
CPU_ROM_MEM[141 ] <= 32'hC00061CC;
CPU_ROM_MEM[142 ] <= 32'hC0006180;
CPU_ROM_MEM[143 ] <= 32'hC0006140;
CPU_ROM_MEM[144 ] <= 32'hC0006100;
CPU_ROM_MEM[145 ] <= 32'hC0006100;
CPU_ROM_MEM[146 ] <= 32'hC0006100;
CPU_ROM_MEM[147 ] <= 32'hC00063FF;
CPU_ROM_MEM[148 ] <= 32'hC00061FF;
CPU_ROM_MEM[149 ] <= 32'hC00061CC;
CPU_ROM_MEM[150 ] <= 32'hC0006180;
CPU_ROM_MEM[151 ] <= 32'hC0006140;
CPU_ROM_MEM[152 ] <= 32'hC0006100;
CPU_ROM_MEM[153 ] <= 32'hC0006100;
CPU_ROM_MEM[154 ] <= 32'hC0006100;
CPU_ROM_MEM[155 ] <= 32'hC00067FF;
CPU_ROM_MEM[156 ] <= 32'hF9BF67FF;
CPU_ROM_MEM[157 ] <= 32'hF9C566FF;
CPU_ROM_MEM[158 ] <= 32'hF9CE66FF;
CPU_ROM_MEM[159 ] <= 32'hF9E300B4;
CPU_ROM_MEM[160 ] <= 32'h00E1A016;
CPU_ROM_MEM[161 ] <= 32'h1EC5000F;
CPU_ROM_MEM[162 ] <= 32'hA0161F1F;
CPU_ROM_MEM[163 ] <= 32'h1EB6A016;
CPU_ROM_MEM[164 ] <= 32'h01951F6A;
CPU_ROM_MEM[165 ] <= 32'hA016013B;
CPU_ROM_MEM[166 ] <= 32'h0096A016;
CPU_ROM_MEM[167 ] <= 32'hC0000087;
CPU_ROM_MEM[168 ] <= 32'h00F0A016;
CPU_ROM_MEM[169 ] <= 32'h1E981FE2;
CPU_ROM_MEM[170 ] <= 32'hA0161F90;
CPU_ROM_MEM[171 ] <= 32'h1E98A016;
CPU_ROM_MEM[172 ] <= 32'h01D81FA6;
CPU_ROM_MEM[173 ] <= 32'hA01600F7;
CPU_ROM_MEM[174 ] <= 32'h00F0A016;
CPU_ROM_MEM[175 ] <= 32'hC0000151;
CPU_ROM_MEM[176 ] <= 32'h0078A016;
CPU_ROM_MEM[177 ] <= 32'h1EDC0087;
CPU_ROM_MEM[178 ] <= 32'hA0161E98;
CPU_ROM_MEM[179 ] <= 32'h1F97A016;
CPU_ROM_MEM[180 ] <= 32'h009E1E7A;
CPU_ROM_MEM[181 ] <= 32'hA01601AB;
CPU_ROM_MEM[182 ] <= 32'h003CA016;
CPU_ROM_MEM[183 ] <= 32'hC0001E82;
CPU_ROM_MEM[184 ] <= 32'h002DA016;
CPU_ROM_MEM[185 ] <= 32'h015100D2;
CPU_ROM_MEM[186 ] <= 32'hA0160151;
CPU_ROM_MEM[187 ] <= 32'h1FA6A016;
CPU_ROM_MEM[188 ] <= 32'h00171ED4;
CPU_ROM_MEM[189 ] <= 32'hA0161EC5;
CPU_ROM_MEM[190 ] <= 32'h1F88A016;
CPU_ROM_MEM[191 ] <= 32'hC000B980;
CPU_ROM_MEM[192 ] <= 32'h45054AE5;
CPU_ROM_MEM[193 ] <= 32'h5BE040E5;
CPU_ROM_MEM[194 ] <= 32'h5BF65B1B;
CPU_ROM_MEM[195 ] <= 32'h5B0556E5;
CPU_ROM_MEM[196 ] <= 32'h45E040E5;
CPU_ROM_MEM[197 ] <= 32'h45F6451B;
CPU_ROM_MEM[198 ] <= 32'h5B1B56FB;
CPU_ROM_MEM[199 ] <= 32'h45E040FB;
CPU_ROM_MEM[200 ] <= 32'h45EA4505;
CPU_ROM_MEM[201 ] <= 32'h451B4AFB;
CPU_ROM_MEM[202 ] <= 32'h5BE040FB;
CPU_ROM_MEM[203 ] <= 32'h5BEA5B05;
CPU_ROM_MEM[204 ] <= 32'h8040C000;
CPU_ROM_MEM[205 ] <= 32'h61800000;
CPU_ROM_MEM[206 ] <= 32'hE000C000;
CPU_ROM_MEM[207 ] <= 32'h80407200;
CPU_ROM_MEM[208 ] <= 32'h61800228;
CPU_ROM_MEM[209 ] <= 32'h01E00000;
CPU_ROM_MEM[210 ] <= 32'hE0001BB0;
CPU_ROM_MEM[211 ] <= 32'h00000000;
CPU_ROM_MEM[212 ] <= 32'hE0000000;
CPU_ROM_MEM[213 ] <= 32'h1C400000;
CPU_ROM_MEM[214 ] <= 32'hE0000450;
CPU_ROM_MEM[215 ] <= 32'h00000000;
CPU_ROM_MEM[216 ] <= 32'hE0008040;
CPU_ROM_MEM[217 ] <= 32'hC0000228;
CPU_ROM_MEM[218 ] <= 32'h01E01BB0;
CPU_ROM_MEM[219 ] <= 32'hE0000000;
CPU_ROM_MEM[220 ] <= 32'hFC400450;
CPU_ROM_MEM[221 ] <= 32'hE0000228;
CPU_ROM_MEM[222 ] <= 32'hE3C08040;
CPU_ROM_MEM[223 ] <= 32'hC0000000;
CPU_ROM_MEM[224 ] <= 32'h1FF940E7;
CPU_ROM_MEM[225 ] <= 32'h00001FF9;
CPU_ROM_MEM[226 ] <= 32'hC0000000;
CPU_ROM_MEM[227 ] <= 32'h1FF940E7;
CPU_ROM_MEM[228 ] <= 32'h00071FF9;
CPU_ROM_MEM[229 ] <= 32'h59E00007;
CPU_ROM_MEM[230 ] <= 32'h0000C000;
CPU_ROM_MEM[231 ] <= 32'h00001FF9;
CPU_ROM_MEM[232 ] <= 32'h0005E002;
CPU_ROM_MEM[233 ] <= 32'h0002E005;
CPU_ROM_MEM[234 ] <= 32'h1FFEE005;
CPU_ROM_MEM[235 ] <= 32'h1FFBE002;
CPU_ROM_MEM[236 ] <= 32'h1FFBFFFE;
CPU_ROM_MEM[237 ] <= 32'h1FFEFFFB;
CPU_ROM_MEM[238 ] <= 32'h0002FFFB;
CPU_ROM_MEM[239 ] <= 32'h0005FFFE;
CPU_ROM_MEM[240 ] <= 32'h00000007;
CPU_ROM_MEM[241 ] <= 32'hC0004019;
CPU_ROM_MEM[242 ] <= 32'h45E242E5;
CPU_ROM_MEM[243 ] <= 32'h5EE55BE2;
CPU_ROM_MEM[244 ] <= 32'h5BFE5EFB;
CPU_ROM_MEM[245 ] <= 32'h42FB45FE;
CPU_ROM_MEM[246 ] <= 32'h4007C000;
CPU_ROM_MEM[247 ] <= 32'hB9EF0000;
CPU_ROM_MEM[248 ] <= 32'hE000C000;
CPU_ROM_MEM[249 ] <= 32'h64800210;
CPU_ROM_MEM[250 ] <= 32'h1E68B88F;
CPU_ROM_MEM[251 ] <= 32'hB841B879;
CPU_ROM_MEM[252 ] <= 32'hB88BB84C;
CPU_ROM_MEM[253 ] <= 32'h80400210;
CPU_ROM_MEM[254 ] <= 32'h0180B8A0;
CPU_ROM_MEM[255 ] <= 32'hB82FB89C;
CPU_ROM_MEM[256 ] <= 32'hB84C8040;
CPU_ROM_MEM[257 ] <= 32'hC00001C8;
CPU_ROM_MEM[258 ] <= 32'h1FB8B88F;
CPU_ROM_MEM[259 ] <= 32'hB85AB85F;
CPU_ROM_MEM[260 ] <= 32'hB84CB86E;
CPU_ROM_MEM[261 ] <= 32'hB8458040;
CPU_ROM_MEM[262 ] <= 32'hC0001F98;
CPU_ROM_MEM[263 ] <= 32'h01E06180;
CPU_ROM_MEM[264 ] <= 32'h001E0064;
CPU_ROM_MEM[265 ] <= 32'h0000FFBA;
CPU_ROM_MEM[266 ] <= 32'h56F60000;
CPU_ROM_MEM[267 ] <= 32'hE05A0000;
CPU_ROM_MEM[268 ] <= 32'h1FA656E0;
CPU_ROM_MEM[269 ] <= 32'h0000E05A;
CPU_ROM_MEM[270 ] <= 32'h00001FA6;
CPU_ROM_MEM[271 ] <= 32'h56EA0000;
CPU_ROM_MEM[272 ] <= 32'hE0466480;
CPU_ROM_MEM[273 ] <= 32'h000A1FB0;
CPU_ROM_MEM[274 ] <= 32'h40F645FB;
CPU_ROM_MEM[275 ] <= 32'h40EA4016;
CPU_ROM_MEM[276 ] <= 32'h4AE040EA;
CPU_ROM_MEM[277 ] <= 32'h401645E5;
CPU_ROM_MEM[278 ] <= 32'h40EA450A;
CPU_ROM_MEM[279 ] <= 32'h4AFB4AF1;
CPU_ROM_MEM[280 ] <= 32'h0000FFC4;
CPU_ROM_MEM[281 ] <= 32'h5BE05BEA;
CPU_ROM_MEM[282 ] <= 32'h56E51FC4;
CPU_ROM_MEM[283 ] <= 32'hE00056FB;
CPU_ROM_MEM[284 ] <= 32'h5BF65BE0;
CPU_ROM_MEM[285 ] <= 32'h0000E03C;
CPU_ROM_MEM[286 ] <= 32'h4AEF4AE5;
CPU_ROM_MEM[287 ] <= 32'h561B0000;
CPU_ROM_MEM[288 ] <= 32'hFFC456F1;
CPU_ROM_MEM[289 ] <= 32'h4A0F4AE5;
CPU_ROM_MEM[290 ] <= 32'h003CE000;
CPU_ROM_MEM[291 ] <= 32'h4AFB0000;
CPU_ROM_MEM[292 ] <= 32'hE03C0000;
CPU_ROM_MEM[293 ] <= 32'h1FC44AF1;
CPU_ROM_MEM[294 ] <= 32'h61801FC4;
CPU_ROM_MEM[295 ] <= 32'h001E0000;
CPU_ROM_MEM[296 ] <= 32'hFFCE5BFB;
CPU_ROM_MEM[297 ] <= 32'h5BE50000;
CPU_ROM_MEM[298 ] <= 32'hE0324500;
CPU_ROM_MEM[299 ] <= 32'h0000FFC4;
CPU_ROM_MEM[300 ] <= 32'h8040C000;
CPU_ROM_MEM[301 ] <= 32'h1DD801E0;
CPU_ROM_MEM[302 ] <= 32'h61801FEC;
CPU_ROM_MEM[303 ] <= 32'h0064001E;
CPU_ROM_MEM[304 ] <= 32'hFFCE40F6;
CPU_ROM_MEM[305 ] <= 32'h56F656E0;
CPU_ROM_MEM[306 ] <= 32'h56EA1FD8;
CPU_ROM_MEM[307 ] <= 32'hE0464500;
CPU_ROM_MEM[308 ] <= 32'h0032FFA6;
CPU_ROM_MEM[309 ] <= 32'h4A001FCE;
CPU_ROM_MEM[310 ] <= 32'hE05A4F00;
CPU_ROM_MEM[311 ] <= 32'h0028FFBA;
CPU_ROM_MEM[312 ] <= 32'h648040F1;
CPU_ROM_MEM[313 ] <= 32'h5BFB56E0;
CPU_ROM_MEM[314 ] <= 32'h5BE55BEA;
CPU_ROM_MEM[315 ] <= 32'h451B45F6;
CPU_ROM_MEM[316 ] <= 32'h4A005BEA;
CPU_ROM_MEM[317 ] <= 32'h450545F6;
CPU_ROM_MEM[318 ] <= 32'h00000028;
CPU_ROM_MEM[319 ] <= 32'h4AE04AFB;
CPU_ROM_MEM[320 ] <= 32'h4AF10000;
CPU_ROM_MEM[321 ] <= 32'hFFC45BE0;
CPU_ROM_MEM[322 ] <= 32'h5BEA56E5;
CPU_ROM_MEM[323 ] <= 32'h1FC4E000;
CPU_ROM_MEM[324 ] <= 32'h56FB5BF6;
CPU_ROM_MEM[325 ] <= 32'h5BE00000;
CPU_ROM_MEM[326 ] <= 32'hE03C4AEF;
CPU_ROM_MEM[327 ] <= 32'h0000FFC4;
CPU_ROM_MEM[328 ] <= 32'h56F14A0F;
CPU_ROM_MEM[329 ] <= 32'h4AE5003C;
CPU_ROM_MEM[330 ] <= 32'hE0004AFB;
CPU_ROM_MEM[331 ] <= 32'h4AF1560F;
CPU_ROM_MEM[332 ] <= 32'h0000E03C;
CPU_ROM_MEM[333 ] <= 32'h61801FE2;
CPU_ROM_MEM[334 ] <= 32'h1FC40014;
CPU_ROM_MEM[335 ] <= 32'hFFD840F6;
CPU_ROM_MEM[336 ] <= 32'h5BE05BE5;
CPU_ROM_MEM[337 ] <= 32'h1FE2E032;
CPU_ROM_MEM[338 ] <= 32'h4500001E;
CPU_ROM_MEM[339 ] <= 32'hFFC44505;
CPU_ROM_MEM[340 ] <= 32'h1FE2E032;
CPU_ROM_MEM[341 ] <= 32'h8040C000;
CPU_ROM_MEM[342 ] <= 32'h1DD80000;
CPU_ROM_MEM[343 ] <= 32'h61801F9C;
CPU_ROM_MEM[344 ] <= 32'h1F88003C;
CPU_ROM_MEM[345 ] <= 32'hE0144AEA;
CPU_ROM_MEM[346 ] <= 32'h4AEF4AEA;
CPU_ROM_MEM[347 ] <= 32'h0000E03C;
CPU_ROM_MEM[348 ] <= 32'h56EA56EF;
CPU_ROM_MEM[349 ] <= 32'h56EA1FC4;
CPU_ROM_MEM[350 ] <= 32'hE0144011;
CPU_ROM_MEM[351 ] <= 32'h003CFFEC;
CPU_ROM_MEM[352 ] <= 32'h0028FFD8;
CPU_ROM_MEM[353 ] <= 32'h0000FFC4;
CPU_ROM_MEM[354 ] <= 32'h1FD8FFD8;
CPU_ROM_MEM[355 ] <= 32'h1FC4FFEC;
CPU_ROM_MEM[356 ] <= 32'h400A6480;
CPU_ROM_MEM[357 ] <= 32'h005AE01E;
CPU_ROM_MEM[358 ] <= 32'h000A0050;
CPU_ROM_MEM[359 ] <= 32'h1F9CE01E;
CPU_ROM_MEM[360 ] <= 32'h00460014;
CPU_ROM_MEM[361 ] <= 32'h4FF60028;
CPU_ROM_MEM[362 ] <= 32'hFFE24AF6;
CPU_ROM_MEM[363 ] <= 32'h1FD8E00A;
CPU_ROM_MEM[364 ] <= 32'h00281FF6;
CPU_ROM_MEM[365 ] <= 32'h0000FFD8;
CPU_ROM_MEM[366 ] <= 32'h1FD8FFF6;
CPU_ROM_MEM[367 ] <= 32'h0028000A;
CPU_ROM_MEM[368 ] <= 32'h56F61FD8;
CPU_ROM_MEM[369 ] <= 32'hFFE251F6;
CPU_ROM_MEM[370 ] <= 32'h8040C000;
CPU_ROM_MEM[371 ] <= 32'h1F981E20;
CPU_ROM_MEM[372 ] <= 32'h6180001E;
CPU_ROM_MEM[373 ] <= 32'h1F9C0000;
CPU_ROM_MEM[374 ] <= 32'hE04656EA;
CPU_ROM_MEM[375 ] <= 32'h0000FFA6;
CPU_ROM_MEM[376 ] <= 32'h0000005A;
CPU_ROM_MEM[377 ] <= 32'h56E00000;
CPU_ROM_MEM[378 ] <= 32'hFFA60000;
CPU_ROM_MEM[379 ] <= 32'h005A56F6;
CPU_ROM_MEM[380 ] <= 32'h0000FFBA;
CPU_ROM_MEM[381 ] <= 32'h6480000A;
CPU_ROM_MEM[382 ] <= 32'h005040EA;
CPU_ROM_MEM[383 ] <= 32'h45E540F6;
CPU_ROM_MEM[384 ] <= 32'h400A4AE0;
CPU_ROM_MEM[385 ] <= 32'h40F6400A;
CPU_ROM_MEM[386 ] <= 32'h45FB40F6;
CPU_ROM_MEM[387 ] <= 32'h45164AE5;
CPU_ROM_MEM[388 ] <= 32'h4AEF0000;
CPU_ROM_MEM[389 ] <= 32'hE03C5BE0;
CPU_ROM_MEM[390 ] <= 32'h5BF656FB;
CPU_ROM_MEM[391 ] <= 32'h1FC4E000;
CPU_ROM_MEM[392 ] <= 32'h56E55BEA;
CPU_ROM_MEM[393 ] <= 32'h5BE00000;
CPU_ROM_MEM[394 ] <= 32'hFFC44AF1;
CPU_ROM_MEM[395 ] <= 32'h4AFB5605;
CPU_ROM_MEM[396 ] <= 32'h0000E03C;
CPU_ROM_MEM[397 ] <= 32'h56EF4A11;
CPU_ROM_MEM[398 ] <= 32'h4AFB003C;
CPU_ROM_MEM[399 ] <= 32'hE0004AE5;
CPU_ROM_MEM[400 ] <= 32'h0000FFC4;
CPU_ROM_MEM[401 ] <= 32'h0000003C;
CPU_ROM_MEM[402 ] <= 32'h4AEF6180;
CPU_ROM_MEM[403 ] <= 32'h1FC41FE2;
CPU_ROM_MEM[404 ] <= 32'h0000E032;
CPU_ROM_MEM[405 ] <= 32'h5BE55BFB;
CPU_ROM_MEM[406 ] <= 32'h0000FFCE;
CPU_ROM_MEM[407 ] <= 32'h45000000;
CPU_ROM_MEM[408 ] <= 32'hE03C8040;
CPU_ROM_MEM[409 ] <= 32'hC0001DD8;
CPU_ROM_MEM[410 ] <= 32'h1E206180;
CPU_ROM_MEM[411 ] <= 32'h1FEC1F9C;
CPU_ROM_MEM[412 ] <= 32'h001EE032;
CPU_ROM_MEM[413 ] <= 32'h40EA56EA;
CPU_ROM_MEM[414 ] <= 32'h56E056F6;
CPU_ROM_MEM[415 ] <= 32'h1FD8FFBA;
CPU_ROM_MEM[416 ] <= 32'h45000032;
CPU_ROM_MEM[417 ] <= 32'hE05A4A00;
CPU_ROM_MEM[418 ] <= 32'h1FCEFFA6;
CPU_ROM_MEM[419 ] <= 32'h4F000028;
CPU_ROM_MEM[420 ] <= 32'hE0466480;
CPU_ROM_MEM[421 ] <= 32'h40EF5BE5;
CPU_ROM_MEM[422 ] <= 32'h56E05BFB;
CPU_ROM_MEM[423 ] <= 32'h5BF64505;
CPU_ROM_MEM[424 ] <= 32'h45EA4A00;
CPU_ROM_MEM[425 ] <= 32'h5BF6451B;
CPU_ROM_MEM[426 ] <= 32'h45EA0000;
CPU_ROM_MEM[427 ] <= 32'h1FD84AE0;
CPU_ROM_MEM[428 ] <= 32'h4AE54AEF;
CPU_ROM_MEM[429 ] <= 32'h0000E03C;
CPU_ROM_MEM[430 ] <= 32'h5BE05BF6;
CPU_ROM_MEM[431 ] <= 32'h56FB1FC4;
CPU_ROM_MEM[432 ] <= 32'hE00056E5;
CPU_ROM_MEM[433 ] <= 32'h5BEA5BE0;
CPU_ROM_MEM[434 ] <= 32'h0000FFC4;
CPU_ROM_MEM[435 ] <= 32'h4AF10000;
CPU_ROM_MEM[436 ] <= 32'hE03C56EF;
CPU_ROM_MEM[437 ] <= 32'h4A114AFB;
CPU_ROM_MEM[438 ] <= 32'h003CE000;
CPU_ROM_MEM[439 ] <= 32'h4AE54AEF;
CPU_ROM_MEM[440 ] <= 32'h56110000;
CPU_ROM_MEM[441 ] <= 32'hFFC46180;
CPU_ROM_MEM[442 ] <= 32'h1FE2003C;
CPU_ROM_MEM[443 ] <= 32'h0014E028;
CPU_ROM_MEM[444 ] <= 32'h40EA5BE0;
CPU_ROM_MEM[445 ] <= 32'h5BFB1FE2;
CPU_ROM_MEM[446 ] <= 32'hFFCE4500;
CPU_ROM_MEM[447 ] <= 32'h001EE03C;
CPU_ROM_MEM[448 ] <= 32'h451B1FE2;
CPU_ROM_MEM[449 ] <= 32'hFFCE8040;
CPU_ROM_MEM[450 ] <= 32'hC0001FD8;
CPU_ROM_MEM[451 ] <= 32'h0000FBAE;
CPU_ROM_MEM[452 ] <= 32'h1FB00000;
CPU_ROM_MEM[453 ] <= 32'hFBAC1F88;
CPU_ROM_MEM[454 ] <= 32'h0000FBAA;
CPU_ROM_MEM[455 ] <= 32'h1F600000;
CPU_ROM_MEM[456 ] <= 32'hFBA81F38;
CPU_ROM_MEM[457 ] <= 32'h0000FBA6;
CPU_ROM_MEM[458 ] <= 32'h1FD80000;
CPU_ROM_MEM[459 ] <= 32'hFBBB1FB0;
CPU_ROM_MEM[460 ] <= 32'h0000FBB9;
CPU_ROM_MEM[461 ] <= 32'h1F880000;
CPU_ROM_MEM[462 ] <= 32'hFBB71F60;
CPU_ROM_MEM[463 ] <= 32'h0000FBB5;
CPU_ROM_MEM[464 ] <= 32'h1F380000;
CPU_ROM_MEM[465 ] <= 32'hFBB31F10;
CPU_ROM_MEM[466 ] <= 32'h0000FBB1;
CPU_ROM_MEM[467 ] <= 32'h00282000;
CPU_ROM_MEM[468 ] <= 32'h00284000;
CPU_ROM_MEM[469 ] <= 32'h00286000;
CPU_ROM_MEM[470 ] <= 32'h00288000;
CPU_ROM_MEM[471 ] <= 32'h0028A000;
CPU_ROM_MEM[472 ] <= 32'hC0000028;
CPU_ROM_MEM[473 ] <= 32'h20000028;
CPU_ROM_MEM[474 ] <= 32'h40000028;
CPU_ROM_MEM[475 ] <= 32'h60000028;
CPU_ROM_MEM[476 ] <= 32'h80000028;
CPU_ROM_MEM[477 ] <= 32'hA0000028;
CPU_ROM_MEM[478 ] <= 32'hC000C000;
CPU_ROM_MEM[479 ] <= 32'hBC0CFCB8;
CPU_ROM_MEM[480 ] <= 32'hBC0DFCB9;
CPU_ROM_MEM[481 ] <= 32'hBC0FFCBB;
CPU_ROM_MEM[482 ] <= 32'hBC11FCBD;
CPU_ROM_MEM[483 ] <= 32'hBC14FCC0;
CPU_ROM_MEM[484 ] <= 32'hBC17FCC3;
CPU_ROM_MEM[485 ] <= 32'hBC1AFCC6;
CPU_ROM_MEM[486 ] <= 32'hBC1DFCC9;
CPU_ROM_MEM[487 ] <= 32'hBC20FCCC;
CPU_ROM_MEM[488 ] <= 32'hBC23FCCF;
CPU_ROM_MEM[489 ] <= 32'hBC26FCD2;
CPU_ROM_MEM[490 ] <= 32'hBC29FCD5;
CPU_ROM_MEM[491 ] <= 32'hBC2CFCD8;
CPU_ROM_MEM[492 ] <= 32'hBC2FFCDB;
CPU_ROM_MEM[493 ] <= 32'hBC32FCDE;
CPU_ROM_MEM[494 ] <= 32'hBC35FCE1;
CPU_ROM_MEM[495 ] <= 32'hBC38FCE4;
CPU_ROM_MEM[496 ] <= 32'hBC3BFCE7;
CPU_ROM_MEM[497 ] <= 32'hBC3EFCEA;
CPU_ROM_MEM[498 ] <= 32'hBC41FCED;
CPU_ROM_MEM[499 ] <= 32'hBC41FCED;
CPU_ROM_MEM[500 ] <= 32'hBC42FCEE;
CPU_ROM_MEM[501 ] <= 32'hBC42FCEE;
CPU_ROM_MEM[502 ] <= 32'hBC45FCF1;
CPU_ROM_MEM[503 ] <= 32'hBC45FCF1;
CPU_ROM_MEM[504 ] <= 32'hBC48FCF4;
CPU_ROM_MEM[505 ] <= 32'hBC48FCF4;
CPU_ROM_MEM[506 ] <= 32'hBC4BFCF7;
CPU_ROM_MEM[507 ] <= 32'hBC4BFCF7;
CPU_ROM_MEM[508 ] <= 32'hBC4EFCFA;
CPU_ROM_MEM[509 ] <= 32'hBC4EFCFA;
CPU_ROM_MEM[510 ] <= 32'hBC51FCFD;
CPU_ROM_MEM[511 ] <= 32'hBC51FCFD;
CPU_ROM_MEM[512 ] <= 32'hBC54FD00;
CPU_ROM_MEM[513 ] <= 32'hBC54FD00;
CPU_ROM_MEM[514 ] <= 32'hBC57FD03;
CPU_ROM_MEM[515 ] <= 32'hBC57FD03;
CPU_ROM_MEM[516 ] <= 32'hBC5AFD06;
CPU_ROM_MEM[517 ] <= 32'hBC5AFD06;
CPU_ROM_MEM[518 ] <= 32'hC000400F;
CPU_ROM_MEM[519 ] <= 32'hFCB6400F;
CPU_ROM_MEM[520 ] <= 32'hFCB20000;
CPU_ROM_MEM[521 ] <= 32'h003CFCB1;
CPU_ROM_MEM[522 ] <= 32'h0000003C;
CPU_ROM_MEM[523 ] <= 32'hFCAD0000;
CPU_ROM_MEM[524 ] <= 32'h005AFCAC;
CPU_ROM_MEM[525 ] <= 32'h0000005A;
CPU_ROM_MEM[526 ] <= 32'hFCA80000;
CPU_ROM_MEM[527 ] <= 32'h0078FCA7;
CPU_ROM_MEM[528 ] <= 32'h00000078;
CPU_ROM_MEM[529 ] <= 32'hFCA30000;
CPU_ROM_MEM[530 ] <= 32'h0096FCA2;
CPU_ROM_MEM[531 ] <= 32'h00000096;
CPU_ROM_MEM[532 ] <= 32'hFC9E0000;
CPU_ROM_MEM[533 ] <= 32'h00B4FC9D;
CPU_ROM_MEM[534 ] <= 32'h000000B4;
CPU_ROM_MEM[535 ] <= 32'hFC990000;
CPU_ROM_MEM[536 ] <= 32'h00D2FC98;
CPU_ROM_MEM[537 ] <= 32'h000000D2;
CPU_ROM_MEM[538 ] <= 32'hFC940000;
CPU_ROM_MEM[539 ] <= 32'h00F0FC93;
CPU_ROM_MEM[540 ] <= 32'h000000F0;
CPU_ROM_MEM[541 ] <= 32'hFC8F0000;
CPU_ROM_MEM[542 ] <= 32'h00F0FC8E;
CPU_ROM_MEM[543 ] <= 32'h000000F0;
CPU_ROM_MEM[544 ] <= 32'hFC8AC000;
CPU_ROM_MEM[545 ] <= 32'h1FF1E01E;
CPU_ROM_MEM[546 ] <= 32'hFC601FE2;
CPU_ROM_MEM[547 ] <= 32'hE03CFC65;
CPU_ROM_MEM[548 ] <= 32'h1FD3E05A;
CPU_ROM_MEM[549 ] <= 32'hFC691FC4;
CPU_ROM_MEM[550 ] <= 32'hE078FC6E;
CPU_ROM_MEM[551 ] <= 32'h1FB5E096;
CPU_ROM_MEM[552 ] <= 32'hFC731FA6;
CPU_ROM_MEM[553 ] <= 32'hE0B4FC78;
CPU_ROM_MEM[554 ] <= 32'h1F97E0D2;
CPU_ROM_MEM[555 ] <= 32'hFC7D1F88;
CPU_ROM_MEM[556 ] <= 32'hE0F0FC82;
CPU_ROM_MEM[557 ] <= 32'h1F79E10E;
CPU_ROM_MEM[558 ] <= 32'hFC87C000;
CPU_ROM_MEM[559 ] <= 32'h1FF1001E;
CPU_ROM_MEM[560 ] <= 32'h000FE000;
CPU_ROM_MEM[561 ] <= 32'hFCB61FE2;
CPU_ROM_MEM[562 ] <= 32'h003C4FE0;
CPU_ROM_MEM[563 ] <= 32'hFCB11FD3;
CPU_ROM_MEM[564 ] <= 32'h005A002D;
CPU_ROM_MEM[565 ] <= 32'hE000FCAC;
CPU_ROM_MEM[566 ] <= 32'h1FC40078;
CPU_ROM_MEM[567 ] <= 32'h003CE000;
CPU_ROM_MEM[568 ] <= 32'hFCA71FB5;
CPU_ROM_MEM[569 ] <= 32'h0096004B;
CPU_ROM_MEM[570 ] <= 32'hE000FCA2;
CPU_ROM_MEM[571 ] <= 32'h1FA600B4;
CPU_ROM_MEM[572 ] <= 32'h005AE000;
CPU_ROM_MEM[573 ] <= 32'hFC9D1F97;
CPU_ROM_MEM[574 ] <= 32'h00D20069;
CPU_ROM_MEM[575 ] <= 32'hE000FC98;
CPU_ROM_MEM[576 ] <= 32'h1F8800F0;
CPU_ROM_MEM[577 ] <= 32'h0078E000;
CPU_ROM_MEM[578 ] <= 32'hFC931F79;
CPU_ROM_MEM[579 ] <= 32'h010E0087;
CPU_ROM_MEM[580 ] <= 32'hE000FC8E;
CPU_ROM_MEM[581 ] <= 32'h1F790000;
CPU_ROM_MEM[582 ] <= 32'h0087E000;
CPU_ROM_MEM[583 ] <= 32'h40F11FF1;
CPU_ROM_MEM[584 ] <= 32'h0000000F;
CPU_ROM_MEM[585 ] <= 32'hE00040F1;
CPU_ROM_MEM[586 ] <= 32'h1FF10000;
CPU_ROM_MEM[587 ] <= 32'h000FE000;
CPU_ROM_MEM[588 ] <= 32'h40F11FA6;
CPU_ROM_MEM[589 ] <= 32'h0000005A;
CPU_ROM_MEM[590 ] <= 32'hE00040F1;
CPU_ROM_MEM[591 ] <= 32'h1FF10000;
CPU_ROM_MEM[592 ] <= 32'h000FE000;
CPU_ROM_MEM[593 ] <= 32'h40F11FF1;
CPU_ROM_MEM[594 ] <= 32'h0000000F;
CPU_ROM_MEM[595 ] <= 32'hE00040F1;
CPU_ROM_MEM[596 ] <= 32'h1FD30000;
CPU_ROM_MEM[597 ] <= 32'h002DE000;
CPU_ROM_MEM[598 ] <= 32'h40F11FF1;
CPU_ROM_MEM[599 ] <= 32'h0000000F;
CPU_ROM_MEM[600 ] <= 32'hE00040F1;
CPU_ROM_MEM[601 ] <= 32'h1FF10000;
CPU_ROM_MEM[602 ] <= 32'h000FE000;
CPU_ROM_MEM[603 ] <= 32'h40F1C000;
CPU_ROM_MEM[604 ] <= 32'hC0004011;
CPU_ROM_MEM[605 ] <= 32'hFD624011;
CPU_ROM_MEM[606 ] <= 32'hFD5E0000;
CPU_ROM_MEM[607 ] <= 32'h1FC4FD5D;
CPU_ROM_MEM[608 ] <= 32'h00001FC4;
CPU_ROM_MEM[609 ] <= 32'hFD590000;
CPU_ROM_MEM[610 ] <= 32'h1FA6FD58;
CPU_ROM_MEM[611 ] <= 32'h00001FA6;
CPU_ROM_MEM[612 ] <= 32'hFD540000;
CPU_ROM_MEM[613 ] <= 32'h1F88FD53;
CPU_ROM_MEM[614 ] <= 32'h00001F88;
CPU_ROM_MEM[615 ] <= 32'hFD4F0000;
CPU_ROM_MEM[616 ] <= 32'h1F6AFD4E;
CPU_ROM_MEM[617 ] <= 32'h00001F6A;
CPU_ROM_MEM[618 ] <= 32'hFD4A0000;
CPU_ROM_MEM[619 ] <= 32'h1F4CFD49;
CPU_ROM_MEM[620 ] <= 32'h00001F4C;
CPU_ROM_MEM[621 ] <= 32'hFD450000;
CPU_ROM_MEM[622 ] <= 32'h1F2EFD44;
CPU_ROM_MEM[623 ] <= 32'h00001F2E;
CPU_ROM_MEM[624 ] <= 32'hFD400000;
CPU_ROM_MEM[625 ] <= 32'h1F10FD3F;
CPU_ROM_MEM[626 ] <= 32'h00001F10;
CPU_ROM_MEM[627 ] <= 32'hFD3B0000;
CPU_ROM_MEM[628 ] <= 32'h1F10FD3A;
CPU_ROM_MEM[629 ] <= 32'h00001F10;
CPU_ROM_MEM[630 ] <= 32'hFD36C000;
CPU_ROM_MEM[631 ] <= 32'h1FF1FFE2;
CPU_ROM_MEM[632 ] <= 32'hFD0C1FE2;
CPU_ROM_MEM[633 ] <= 32'hFFC4FD11;
CPU_ROM_MEM[634 ] <= 32'h1FD3FFA6;
CPU_ROM_MEM[635 ] <= 32'hFD151FC4;
CPU_ROM_MEM[636 ] <= 32'hFF88FD1A;
CPU_ROM_MEM[637 ] <= 32'h1FB5FF6A;
CPU_ROM_MEM[638 ] <= 32'hFD1F1FA6;
CPU_ROM_MEM[639 ] <= 32'hFF4CFD24;
CPU_ROM_MEM[640 ] <= 32'h1F97FF2E;
CPU_ROM_MEM[641 ] <= 32'hFD291F88;
CPU_ROM_MEM[642 ] <= 32'hFF10FD2E;
CPU_ROM_MEM[643 ] <= 32'h1F79FEF2;
CPU_ROM_MEM[644 ] <= 32'hFD33C000;
CPU_ROM_MEM[645 ] <= 32'h1FF11FE2;
CPU_ROM_MEM[646 ] <= 32'h000FE000;
CPU_ROM_MEM[647 ] <= 32'hFD621FE2;
CPU_ROM_MEM[648 ] <= 32'h1FC44FE0;
CPU_ROM_MEM[649 ] <= 32'hFD5D1FD3;
CPU_ROM_MEM[650 ] <= 32'h1FA6002D;
CPU_ROM_MEM[651 ] <= 32'hE000FD58;
CPU_ROM_MEM[652 ] <= 32'h1FC41F88;
CPU_ROM_MEM[653 ] <= 32'h003CE000;
CPU_ROM_MEM[654 ] <= 32'hFD531FB5;
CPU_ROM_MEM[655 ] <= 32'h1F6A004B;
CPU_ROM_MEM[656 ] <= 32'hE000FD4E;
CPU_ROM_MEM[657 ] <= 32'h1FA61F4C;
CPU_ROM_MEM[658 ] <= 32'h005AE000;
CPU_ROM_MEM[659 ] <= 32'hFD491F97;
CPU_ROM_MEM[660 ] <= 32'h1F2E0069;
CPU_ROM_MEM[661 ] <= 32'hE000FD44;
CPU_ROM_MEM[662 ] <= 32'h1F881F10;
CPU_ROM_MEM[663 ] <= 32'h0078E000;
CPU_ROM_MEM[664 ] <= 32'hFD3F1F79;
CPU_ROM_MEM[665 ] <= 32'h1EF20087;
CPU_ROM_MEM[666 ] <= 32'hE000FD3A;
CPU_ROM_MEM[667 ] <= 32'h1F790000;
CPU_ROM_MEM[668 ] <= 32'h0087E000;
CPU_ROM_MEM[669 ] <= 32'h40EF1FF1;
CPU_ROM_MEM[670 ] <= 32'h0000000F;
CPU_ROM_MEM[671 ] <= 32'hE00040EF;
CPU_ROM_MEM[672 ] <= 32'h1FF10000;
CPU_ROM_MEM[673 ] <= 32'h000FE000;
CPU_ROM_MEM[674 ] <= 32'h40EF1FA6;
CPU_ROM_MEM[675 ] <= 32'h0000005A;
CPU_ROM_MEM[676 ] <= 32'hE00040EF;
CPU_ROM_MEM[677 ] <= 32'h1FF10000;
CPU_ROM_MEM[678 ] <= 32'h000FE000;
CPU_ROM_MEM[679 ] <= 32'h40EF1FF1;
CPU_ROM_MEM[680 ] <= 32'h0000000F;
CPU_ROM_MEM[681 ] <= 32'hE00040EF;
CPU_ROM_MEM[682 ] <= 32'h1FD30000;
CPU_ROM_MEM[683 ] <= 32'h002DE000;
CPU_ROM_MEM[684 ] <= 32'h40EF1FF1;
CPU_ROM_MEM[685 ] <= 32'h0000000F;
CPU_ROM_MEM[686 ] <= 32'hE00040EF;
CPU_ROM_MEM[687 ] <= 32'h1FF10000;
CPU_ROM_MEM[688 ] <= 32'h000FE000;
CPU_ROM_MEM[689 ] <= 32'h40EFC000;
CPU_ROM_MEM[690 ] <= 32'h62801E20;
CPU_ROM_MEM[691 ] <= 32'h0620FD83;
CPU_ROM_MEM[692 ] <= 32'h62801E20;
CPU_ROM_MEM[693 ] <= 32'h19E01E20;
CPU_ROM_MEM[694 ] <= 32'hA0601E20;
CPU_ROM_MEM[695 ] <= 32'hA0C01E20;
CPU_ROM_MEM[696 ] <= 32'hA1401EE0;
CPU_ROM_MEM[697 ] <= 32'hA1401F70;
CPU_ROM_MEM[698 ] <= 32'hA1401FD0;
CPU_ROM_MEM[699 ] <= 32'hA1400030;
CPU_ROM_MEM[700 ] <= 32'hA1400090;
CPU_ROM_MEM[701 ] <= 32'hA1400120;
CPU_ROM_MEM[702 ] <= 32'hA14001E0;
CPU_ROM_MEM[703 ] <= 32'hA14001E0;
CPU_ROM_MEM[704 ] <= 32'hC0C001E0;
CPU_ROM_MEM[705 ] <= 32'hC06001E0;
CPU_ROM_MEM[706 ] <= 32'hE02001E0;
CPU_ROM_MEM[707 ] <= 32'hFFE001E0;
CPU_ROM_MEM[708 ] <= 32'hFFA001E0;
CPU_ROM_MEM[709 ] <= 32'hFF4001E0;
CPU_ROM_MEM[710 ] <= 32'hFEC00120;
CPU_ROM_MEM[711 ] <= 32'hFEC00090;
CPU_ROM_MEM[712 ] <= 32'hDEC00030;
CPU_ROM_MEM[713 ] <= 32'hDEC01FD0;
CPU_ROM_MEM[714 ] <= 32'hBEC01F70;
CPU_ROM_MEM[715 ] <= 32'hBEC01EE0;
CPU_ROM_MEM[716 ] <= 32'hBEC01E20;
CPU_ROM_MEM[717 ] <= 32'hBEC01E20;
CPU_ROM_MEM[718 ] <= 32'hBF401E20;
CPU_ROM_MEM[719 ] <= 32'hBFA01E20;
CPU_ROM_MEM[720 ] <= 32'hBFE01E20;
CPU_ROM_MEM[721 ] <= 32'hA0207200;
CPU_ROM_MEM[722 ] <= 32'h8040C000;
CPU_ROM_MEM[723 ] <= 32'h678001E0;
CPU_ROM_MEM[724 ] <= 32'h06201C70;
CPU_ROM_MEM[725 ] <= 32'hD3C01FD0;
CPU_ROM_MEM[726 ] <= 32'h00000390;
CPU_ROM_MEM[727 ] <= 32'hCC407200;
CPU_ROM_MEM[728 ] <= 32'h8040C000;
CPU_ROM_MEM[729 ] <= 32'h64800330;
CPU_ROM_MEM[730 ] <= 32'h02800060;
CPU_ROM_MEM[731 ] <= 32'hDF800090;
CPU_ROM_MEM[732 ] <= 32'hDFA000C0;
CPU_ROM_MEM[733 ] <= 32'hDFC000C0;
CPU_ROM_MEM[734 ] <= 32'hDFE000C0;
CPU_ROM_MEM[735 ] <= 32'hC0200090;
CPU_ROM_MEM[736 ] <= 32'hC0600030;
CPU_ROM_MEM[737 ] <= 32'hC0800000;
CPU_ROM_MEM[738 ] <= 32'hC0801FA0;
CPU_ROM_MEM[739 ] <= 32'hC0801F40;
CPU_ROM_MEM[740 ] <= 32'hC0801F40;
CPU_ROM_MEM[741 ] <= 32'hC0601F40;
CPU_ROM_MEM[742 ] <= 32'hC0201F40;
CPU_ROM_MEM[743 ] <= 32'hDFE01F70;
CPU_ROM_MEM[744 ] <= 32'hDFA01FD0;
CPU_ROM_MEM[745 ] <= 32'hDF800000;
CPU_ROM_MEM[746 ] <= 32'hDFA00030;
CPU_ROM_MEM[747 ] <= 32'hDFA07200;
CPU_ROM_MEM[748 ] <= 32'h8040C000;
CPU_ROM_MEM[749 ] <= 32'h64800330;
CPU_ROM_MEM[750 ] <= 32'h028001E0;
CPU_ROM_MEM[751 ] <= 32'hA0401E80;
CPU_ROM_MEM[752 ] <= 32'hBF400090;
CPU_ROM_MEM[753 ] <= 32'h1FA000F0;
CPU_ROM_MEM[754 ] <= 32'hA1201FD0;
CPU_ROM_MEM[755 ] <= 32'hBEA000C0;
CPU_ROM_MEM[756 ] <= 32'h1FE01F70;
CPU_ROM_MEM[757 ] <= 32'hA1800150;
CPU_ROM_MEM[758 ] <= 32'hBEA00090;
CPU_ROM_MEM[759 ] <= 32'h00601E20;
CPU_ROM_MEM[760 ] <= 32'hA1000210;
CPU_ROM_MEM[761 ] <= 32'hBF800000;
CPU_ROM_MEM[762 ] <= 32'h00801DF0;
CPU_ROM_MEM[763 ] <= 32'hA00001B0;
CPU_ROM_MEM[764 ] <= 32'hA0801C70;
CPU_ROM_MEM[765 ] <= 32'h008001E0;
CPU_ROM_MEM[766 ] <= 32'hBF001DF0;
CPU_ROM_MEM[767 ] <= 32'hA0800000;
CPU_ROM_MEM[768 ] <= 32'h1FA00210;
CPU_ROM_MEM[769 ] <= 32'hBFE07200;
CPU_ROM_MEM[770 ] <= 32'h8040C000;
CPU_ROM_MEM[771 ] <= 32'h628008D0;
CPU_ROM_MEM[772 ] <= 32'h01E01F40;
CPU_ROM_MEM[773 ] <= 32'hA0400030;
CPU_ROM_MEM[774 ] <= 32'hA0800030;
CPU_ROM_MEM[775 ] <= 32'h00001EB0;
CPU_ROM_MEM[776 ] <= 32'hA0600060;
CPU_ROM_MEM[777 ] <= 32'h1FE00030;
CPU_ROM_MEM[778 ] <= 32'hA0801E80;
CPU_ROM_MEM[779 ] <= 32'hA06000C0;
CPU_ROM_MEM[780 ] <= 32'h00401AF0;
CPU_ROM_MEM[781 ] <= 32'hA1800030;
CPU_ROM_MEM[782 ] <= 32'hA0800390;
CPU_ROM_MEM[783 ] <= 32'hBEE01DF0;
CPU_ROM_MEM[784 ] <= 32'h00201FD0;
CPU_ROM_MEM[785 ] <= 32'hBF8000F0;
CPU_ROM_MEM[786 ] <= 32'h1FC01E20;
CPU_ROM_MEM[787 ] <= 32'hA0801FD0;
CPU_ROM_MEM[788 ] <= 32'hBF8000F0;
CPU_ROM_MEM[789 ] <= 32'hBFC01F10;
CPU_ROM_MEM[790 ] <= 32'h00401FD0;
CPU_ROM_MEM[791 ] <= 32'hBF8000F0;
CPU_ROM_MEM[792 ] <= 32'hBFC01C10;
CPU_ROM_MEM[793 ] <= 32'h01400150;
CPU_ROM_MEM[794 ] <= 32'hBFC00030;
CPU_ROM_MEM[795 ] <= 32'hA0800030;
CPU_ROM_MEM[796 ] <= 32'h00800030;
CPU_ROM_MEM[797 ] <= 32'hA0801EE0;
CPU_ROM_MEM[798 ] <= 32'hA0401E20;
CPU_ROM_MEM[799 ] <= 32'h1FC00360;
CPU_ROM_MEM[800 ] <= 32'hBF601FD0;
CPU_ROM_MEM[801 ] <= 32'hBF801B80;
CPU_ROM_MEM[802 ] <= 32'hA0E000F0;
CPU_ROM_MEM[803 ] <= 32'h00401FD0;
CPU_ROM_MEM[804 ] <= 32'hBFA000F0;
CPU_ROM_MEM[805 ] <= 32'h1F600030;
CPU_ROM_MEM[806 ] <= 32'hA0607200;
CPU_ROM_MEM[807 ] <= 32'h8040C000;
CPU_ROM_MEM[808 ] <= 32'h6780000F;
CPU_ROM_MEM[809 ] <= 32'h00311FE2;
CPU_ROM_MEM[810 ] <= 32'hDF9E6280;
CPU_ROM_MEM[811 ] <= 32'h1FE2A009;
CPU_ROM_MEM[812 ] <= 32'h54AA5DAA;
CPU_ROM_MEM[813 ] <= 32'h43AA4CAA;
CPU_ROM_MEM[814 ] <= 32'h001EC009;
CPU_ROM_MEM[815 ] <= 32'h4FE0001E;
CPU_ROM_MEM[816 ] <= 32'hFFF74CF6;
CPU_ROM_MEM[817 ] <= 32'h43D65DB6;
CPU_ROM_MEM[818 ] <= 32'h54B61FE2;
CPU_ROM_MEM[819 ] <= 32'hBFF751A0;
CPU_ROM_MEM[820 ] <= 32'h6480002D;
CPU_ROM_MEM[821 ] <= 32'h00521FFA;
CPU_ROM_MEM[822 ] <= 32'hDFF90001;
CPU_ROM_MEM[823 ] <= 32'hDFFA0008;
CPU_ROM_MEM[824 ] <= 32'hDFF9000C;
CPU_ROM_MEM[825 ] <= 32'hDFFD45C2;
CPU_ROM_MEM[826 ] <= 32'h41C41FF1;
CPU_ROM_MEM[827 ] <= 32'hC00B5AC0;
CPU_ROM_MEM[828 ] <= 32'h64800015;
CPU_ROM_MEM[829 ] <= 32'hBFEA0006;
CPU_ROM_MEM[830 ] <= 32'h000B50A0;
CPU_ROM_MEM[831 ] <= 32'h00081FF7;
CPU_ROM_MEM[832 ] <= 32'h0007A009;
CPU_ROM_MEM[833 ] <= 32'h62800018;
CPU_ROM_MEM[834 ] <= 32'h1FFB1FF7;
CPU_ROM_MEM[835 ] <= 32'hA00F1FE5;
CPU_ROM_MEM[836 ] <= 32'hA0085ABB;
CPU_ROM_MEM[837 ] <= 32'h5A051FE1;
CPU_ROM_MEM[838 ] <= 32'hA0067200;
CPU_ROM_MEM[839 ] <= 32'h8040C000;
CPU_ROM_MEM[840 ] <= 32'h00004100;
CPU_ROM_MEM[841 ] <= 32'h00101F00;
CPU_ROM_MEM[842 ] <= 32'h00006100;
CPU_ROM_MEM[843 ] <= 32'h00101F00;
CPU_ROM_MEM[844 ] <= 32'h00008100;
CPU_ROM_MEM[845 ] <= 32'h00101F00;
CPU_ROM_MEM[846 ] <= 32'h0000A100;
CPU_ROM_MEM[847 ] <= 32'h00101F00;
CPU_ROM_MEM[848 ] <= 32'h0000C100;
CPU_ROM_MEM[849 ] <= 32'h00101F00;
CPU_ROM_MEM[850 ] <= 32'h0000E100;
CPU_ROM_MEM[851 ] <= 32'hC000BFAE;
CPU_ROM_MEM[852 ] <= 32'h80400040;
CPU_ROM_MEM[853 ] <= 32'h1E806480;
CPU_ROM_MEM[854 ] <= 32'hBE908040;
CPU_ROM_MEM[855 ] <= 32'h00401F80;
CPU_ROM_MEM[856 ] <= 32'h6180BE90;
CPU_ROM_MEM[857 ] <= 32'h80400040;
CPU_ROM_MEM[858 ] <= 32'h00806280;
CPU_ROM_MEM[859 ] <= 32'hBE908040;
CPU_ROM_MEM[860 ] <= 32'h1F601E80;
CPU_ROM_MEM[861 ] <= 32'h6680BE90;
CPU_ROM_MEM[862 ] <= 32'h80401F60;
CPU_ROM_MEM[863 ] <= 32'h1F806380;
CPU_ROM_MEM[864 ] <= 32'hBE908040;
CPU_ROM_MEM[865 ] <= 32'h1F600080;
CPU_ROM_MEM[866 ] <= 32'h6580BE90;
CPU_ROM_MEM[867 ] <= 32'h80401FD0;
CPU_ROM_MEM[868 ] <= 32'h1F806780;
CPU_ROM_MEM[869 ] <= 32'hBE908040;
CPU_ROM_MEM[870 ] <= 32'h1F400080;
CPU_ROM_MEM[871 ] <= 32'h67000000;
CPU_ROM_MEM[872 ] <= 32'hE1001FEC;
CPU_ROM_MEM[873 ] <= 32'h1F006710;
CPU_ROM_MEM[874 ] <= 32'h0000E100;
CPU_ROM_MEM[875 ] <= 32'h1FEC1F00;
CPU_ROM_MEM[876 ] <= 32'h67200000;
CPU_ROM_MEM[877 ] <= 32'hE1001FEC;
CPU_ROM_MEM[878 ] <= 32'h1F006730;
CPU_ROM_MEM[879 ] <= 32'h0000E100;
CPU_ROM_MEM[880 ] <= 32'h1FEC1F00;
CPU_ROM_MEM[881 ] <= 32'h67400000;
CPU_ROM_MEM[882 ] <= 32'hE1001FEC;
CPU_ROM_MEM[883 ] <= 32'h1F006750;
CPU_ROM_MEM[884 ] <= 32'h0000E100;
CPU_ROM_MEM[885 ] <= 32'h1FEC1F00;
CPU_ROM_MEM[886 ] <= 32'h67600000;
CPU_ROM_MEM[887 ] <= 32'hE1001FEC;
CPU_ROM_MEM[888 ] <= 32'h1F006770;
CPU_ROM_MEM[889 ] <= 32'h0000E100;
CPU_ROM_MEM[890 ] <= 32'h1FEC1F00;
CPU_ROM_MEM[891 ] <= 32'h67800000;
CPU_ROM_MEM[892 ] <= 32'hE1001FEC;
CPU_ROM_MEM[893 ] <= 32'h1F008040;
CPU_ROM_MEM[894 ] <= 32'hC000BFAE;
CPU_ROM_MEM[895 ] <= 32'h80401DD8;
CPU_ROM_MEM[896 ] <= 32'h1E200450;
CPU_ROM_MEM[897 ] <= 32'hE2D01E90;
CPU_ROM_MEM[898 ] <= 32'hE0F01D20;
CPU_ROM_MEM[899 ] <= 32'hFE2002E0;
CPU_ROM_MEM[900 ] <= 32'hFE200170;
CPU_ROM_MEM[901 ] <= 32'hE0F01BB0;
CPU_ROM_MEM[902 ] <= 32'hE2D00450;
CPU_ROM_MEM[903 ] <= 32'h00001BB0;
CPU_ROM_MEM[904 ] <= 32'hFD300170;
CPU_ROM_MEM[905 ] <= 32'hFF1002E0;
CPU_ROM_MEM[906 ] <= 32'hE1E01D20;
CPU_ROM_MEM[907 ] <= 32'hE1E01E90;
CPU_ROM_MEM[908 ] <= 32'hFF100450;
CPU_ROM_MEM[909 ] <= 32'hFD308040;
CPU_ROM_MEM[910 ] <= 32'h1E9A1E20;
CPU_ROM_MEM[911 ] <= 32'h7240F801;
CPU_ROM_MEM[912 ] <= 32'h72008040;
CPU_ROM_MEM[913 ] <= 32'h1DF101E0;
CPU_ROM_MEM[914 ] <= 32'h0000FC40;
CPU_ROM_MEM[915 ] <= 32'h80401E51;
CPU_ROM_MEM[916 ] <= 32'h01E00000;
CPU_ROM_MEM[917 ] <= 32'hFC408040;
CPU_ROM_MEM[918 ] <= 32'h1EB101E0;
CPU_ROM_MEM[919 ] <= 32'h0000FC40;
CPU_ROM_MEM[920 ] <= 32'h80401F11;
CPU_ROM_MEM[921 ] <= 32'h01E00000;
CPU_ROM_MEM[922 ] <= 32'hFC408040;
CPU_ROM_MEM[923 ] <= 32'h1F7101E0;
CPU_ROM_MEM[924 ] <= 32'h0000FC40;
CPU_ROM_MEM[925 ] <= 32'h80401FD1;
CPU_ROM_MEM[926 ] <= 32'h01E00000;
CPU_ROM_MEM[927 ] <= 32'hFC408040;
CPU_ROM_MEM[928 ] <= 32'h003101E0;
CPU_ROM_MEM[929 ] <= 32'h0000FC40;
CPU_ROM_MEM[930 ] <= 32'h80400091;
CPU_ROM_MEM[931 ] <= 32'h01E00000;
CPU_ROM_MEM[932 ] <= 32'hFC408040;
CPU_ROM_MEM[933 ] <= 32'h00F101E0;
CPU_ROM_MEM[934 ] <= 32'h0000FC40;
CPU_ROM_MEM[935 ] <= 32'h80400151;
CPU_ROM_MEM[936 ] <= 32'h01E00000;
CPU_ROM_MEM[937 ] <= 32'hFC408040;
CPU_ROM_MEM[938 ] <= 32'h01B101E0;
CPU_ROM_MEM[939 ] <= 32'h0000FC40;
CPU_ROM_MEM[940 ] <= 32'h80400211;
CPU_ROM_MEM[941 ] <= 32'h01E00000;
CPU_ROM_MEM[942 ] <= 32'hFC408040;
CPU_ROM_MEM[943 ] <= 32'h02101E21;
CPU_ROM_MEM[944 ] <= 32'h1BE0E000;
CPU_ROM_MEM[945 ] <= 32'h80400210;
CPU_ROM_MEM[946 ] <= 32'h1E611BE0;
CPU_ROM_MEM[947 ] <= 32'hE0008040;
CPU_ROM_MEM[948 ] <= 32'h02101EA1;
CPU_ROM_MEM[949 ] <= 32'h1BE0E000;
CPU_ROM_MEM[950 ] <= 32'h80400210;
CPU_ROM_MEM[951 ] <= 32'h1EE11BE0;
CPU_ROM_MEM[952 ] <= 32'hE0008040;
CPU_ROM_MEM[953 ] <= 32'h02101F21;
CPU_ROM_MEM[954 ] <= 32'h1BE0E000;
CPU_ROM_MEM[955 ] <= 32'h80400210;
CPU_ROM_MEM[956 ] <= 32'h1F611BE0;
CPU_ROM_MEM[957 ] <= 32'hE0008040;
CPU_ROM_MEM[958 ] <= 32'h02101FA1;
CPU_ROM_MEM[959 ] <= 32'h1BE0E000;
CPU_ROM_MEM[960 ] <= 32'h80400210;
CPU_ROM_MEM[961 ] <= 32'h1FE11BE0;
CPU_ROM_MEM[962 ] <= 32'hE0008040;
CPU_ROM_MEM[963 ] <= 32'h02100021;
CPU_ROM_MEM[964 ] <= 32'h1BE0E000;
CPU_ROM_MEM[965 ] <= 32'h80400210;
CPU_ROM_MEM[966 ] <= 32'h00611BE0;
CPU_ROM_MEM[967 ] <= 32'hE0008040;
CPU_ROM_MEM[968 ] <= 32'h021000A1;
CPU_ROM_MEM[969 ] <= 32'h1BE0E000;
CPU_ROM_MEM[970 ] <= 32'h80400210;
CPU_ROM_MEM[971 ] <= 32'h00E11BE0;
CPU_ROM_MEM[972 ] <= 32'hE0008040;
CPU_ROM_MEM[973 ] <= 32'h02100121;
CPU_ROM_MEM[974 ] <= 32'h1BE0E000;
CPU_ROM_MEM[975 ] <= 32'h80400210;
CPU_ROM_MEM[976 ] <= 32'h01611BE0;
CPU_ROM_MEM[977 ] <= 32'hE0008040;
CPU_ROM_MEM[978 ] <= 32'h021001A1;
CPU_ROM_MEM[979 ] <= 32'h1BE0E000;
CPU_ROM_MEM[980 ] <= 32'h80400210;
CPU_ROM_MEM[981 ] <= 32'h01E11BE0;
CPU_ROM_MEM[982 ] <= 32'hE000C000;
CPU_ROM_MEM[983 ] <= 32'h62507200;
CPU_ROM_MEM[984 ] <= 32'h80401DD8;
CPU_ROM_MEM[985 ] <= 32'h1E200000;
CPU_ROM_MEM[986 ] <= 32'hE3C00450;
CPU_ROM_MEM[987 ] <= 32'hE0000000;
CPU_ROM_MEM[988 ] <= 32'hFC401BB0;
CPU_ROM_MEM[989 ] <= 32'hE000C000;
CPU_ROM_MEM[990 ] <= 32'h008A005C;
CPU_ROM_MEM[991 ] <= 32'h0000FF48;
CPU_ROM_MEM[992 ] <= 32'h1EECE000;
CPU_ROM_MEM[993 ] <= 32'h0000E0B8;
CPU_ROM_MEM[994 ] <= 32'h0114E000;
CPU_ROM_MEM[995 ] <= 32'h8040C000;
CPU_ROM_MEM[996 ] <= 32'hBFAF8040;
CPU_ROM_MEM[997 ] <= 32'h01001E20;
CPU_ROM_MEM[998 ] <= 32'h0000E3C0;
CPU_ROM_MEM[999 ] <= 32'h1FFB0000;
CPU_ROM_MEM[1000] <= 32'h0000FC40;
CPU_ROM_MEM[1001] <= 32'h1FFB0000;
CPU_ROM_MEM[1002] <= 32'hC000000C;
CPU_ROM_MEM[1003] <= 32'h01386480;
CPU_ROM_MEM[1004] <= 32'h54E040E8;
CPU_ROM_MEM[1005] <= 32'h4CE040F8;
CPU_ROM_MEM[1006] <= 32'h6280006C;
CPU_ROM_MEM[1007] <= 32'h1FA81F10;
CPU_ROM_MEM[1008] <= 32'hE0005408;
CPU_ROM_MEM[1009] <= 32'h0000E0A0;
CPU_ROM_MEM[1010] <= 32'h4C0800F0;
CPU_ROM_MEM[1011] <= 32'hE0004C18;
CPU_ROM_MEM[1012] <= 32'h0000FF60;
CPU_ROM_MEM[1013] <= 32'h67800030;
CPU_ROM_MEM[1014] <= 32'h1FD01E80;
CPU_ROM_MEM[1015] <= 32'hE0000000;
CPU_ROM_MEM[1016] <= 32'hE1000180;
CPU_ROM_MEM[1017] <= 32'hE0000000;
CPU_ROM_MEM[1018] <= 32'hFF008040;
CPU_ROM_MEM[1019] <= 32'hC0000000;
CPU_ROM_MEM[1020] <= 32'h00000000;
CPU_ROM_MEM[1021] <= 32'h00000000;
CPU_ROM_MEM[1022] <= 32'h00000000;
CPU_ROM_MEM[1023] <= 32'h00000000;
end

reg [31:0] q_a_reg;
always @(posedge clk_a) begin
    q_a_reg <= CPU_ROM_MEM[address_a[11:2]];
end

always @* begin
	case (address_a[1:0]) 
		2'b00 : q_a <= q_a_reg[31:24];
		2'b01 : q_a <= q_a_reg[23:16];
		2'b10 : q_a <= q_a_reg[15:8];
		2'b11 : q_a <= q_a_reg[7:0];
	endcase
end

always @(posedge clk_b) begin
	if (write_b && mask_b[3]) CPU_ROM_MEM[address_b] <= data_b[31:24];
	if (write_b && mask_b[2]) CPU_ROM_MEM[address_b] <= data_b[23:16];
	if (write_b && mask_b[1]) CPU_ROM_MEM[address_b] <= data_b[15:8];
	if (write_b && mask_b[0]) CPU_ROM_MEM[address_b] <= data_b[7:0] ;
	q_b <= CPU_ROM_MEM[address_b];
end

    
endmodule
